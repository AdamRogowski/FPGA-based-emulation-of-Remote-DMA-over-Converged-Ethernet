-- https://docs.amd.com/r/en-US/ug901-vivado-synthesis/Dual-Port-Block-RAM-with-Two-Write-Ports-in-Read-First-Mode-VHDL

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity bram_model is
  generic (
    DATA_WIDTH : integer := 128;
    ADDR_WIDTH : integer := 18; -- 262k locations
    LATENCY    : integer := 3   -- number of pipeline stages
  );
  port (
    clk   : in  std_logic;
    ena   : in  std_logic;
    enb   : in  std_logic;
    wea   : in  std_logic;
    web   : in  std_logic;
    addra : in  std_logic_vector(ADDR_WIDTH - 1 downto 0);
    addrb : in  std_logic_vector(ADDR_WIDTH - 1 downto 0);
    dia   : in  std_logic_vector(DATA_WIDTH - 1 downto 0);
    dib   : in  std_logic_vector(DATA_WIDTH - 1 downto 0);
    doa   : out std_logic_vector(DATA_WIDTH - 1 downto 0);
    dob   : out std_logic_vector(DATA_WIDTH - 1 downto 0)
  );
end entity;

architecture rtl of bram_model is

  -- Memory
  type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(DATA_WIDTH - 1 downto 0);

  constant INIT_BRAM : ram_type := (
    0   => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    1   => "10000000000000000000000000000000000110010000000000011001000000000010000000000000000000000001",
    2   => "10000000000000000000010100000000000110010000000000011001000000000011000000000000000000000010",
    3   => "10000000000000000000101000000000000110010000000000011001000000000100000000000000000000000011",
    4   => "10000000000000000000111100000000000110010000000000011001000111111111000000000000000000000100",
    5   => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    6   => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    7   => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    8   => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    9   => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    10  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    11  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    12  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    13  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    14  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    15  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    16  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    17  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    18  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    19  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    20  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    21  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    22  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    23  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    24  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    25  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    26  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    27  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    28  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    29  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    30  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    31  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    32  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    33  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    34  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    35  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    36  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    37  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    38  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    39  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    40  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    41  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    42  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    43  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    44  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    45  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    46  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    47  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    48  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    49  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    50  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    51  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    52  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    53  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    54  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    55  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    56  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    57  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    58  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    59  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    60  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    61  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    62  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    63  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    64  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    65  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    66  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    67  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    68  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    69  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    70  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    71  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    72  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    73  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    74  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    75  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    76  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    77  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    78  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    79  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    80  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    81  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    82  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    83  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    84  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    85  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    86  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    87  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    88  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    89  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    90  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    91  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    92  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    93  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    94  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    95  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    96  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    97  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    98  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    99  => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    100 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    101 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    102 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    103 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    104 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    105 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    106 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    107 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    108 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    109 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    110 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    111 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    112 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    113 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    114 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    115 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    116 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    117 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    118 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    119 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    120 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    121 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    122 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    123 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    124 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    125 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    126 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    127 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    128 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    129 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    130 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    131 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    132 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    133 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    134 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    135 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    136 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    137 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    138 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    139 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    140 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    141 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    142 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    143 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    144 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    145 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    146 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    147 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    148 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    149 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    150 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    151 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    152 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    153 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    154 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    155 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    156 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    157 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    158 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    159 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    160 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    161 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    162 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    163 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    164 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    165 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    166 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    167 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    168 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    169 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    170 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    171 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    172 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    173 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    174 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    175 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    176 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    177 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    178 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    179 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    180 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    181 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    182 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    183 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    184 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    185 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    186 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    187 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    188 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    189 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    190 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    191 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    192 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    193 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    194 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    195 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    196 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    197 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    198 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    199 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    200 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    201 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    202 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    203 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    204 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    205 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    206 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    207 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    208 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    209 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    210 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    211 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    212 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    213 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    214 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    215 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    216 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    217 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    218 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    219 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    220 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    221 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    222 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    223 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    224 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    225 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    226 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    227 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    228 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    229 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    230 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    231 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    232 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    233 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    234 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    235 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    236 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    237 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    238 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    239 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    240 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    241 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    242 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    243 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    244 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    245 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    246 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    247 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    248 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    249 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    250 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    251 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    252 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    253 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    254 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    255 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    256 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    257 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    258 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    259 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    260 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    261 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    262 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    263 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    264 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    265 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    266 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    267 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    268 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    269 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    270 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    271 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    272 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    273 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    274 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    275 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    276 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    277 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    278 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    279 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    280 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    281 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    282 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    283 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    284 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    285 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    286 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    287 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    288 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    289 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    290 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    291 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    292 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    293 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    294 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    295 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    296 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    297 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    298 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    299 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    300 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    301 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    302 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    303 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    304 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    305 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    306 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    307 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    308 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    309 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    310 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    311 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    312 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    313 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    314 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    315 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    316 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    317 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    318 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    319 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    320 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    321 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    322 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    323 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    324 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    325 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    326 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    327 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    328 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    329 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    330 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    331 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    332 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    333 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    334 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    335 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    336 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    337 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    338 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    339 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    340 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    341 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    342 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    343 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    344 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    345 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    346 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    347 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    348 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    349 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    350 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    351 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    352 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    353 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    354 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    355 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    356 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    357 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    358 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    359 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    360 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    361 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    362 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    363 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    364 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    365 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    366 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    367 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    368 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    369 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    370 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    371 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    372 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    373 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    374 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    375 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    376 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    377 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    378 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    379 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    380 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    381 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    382 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    383 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    384 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    385 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    386 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    387 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    388 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    389 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    390 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    391 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    392 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    393 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    394 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    395 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    396 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    397 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    398 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    399 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    400 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    401 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    402 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    403 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    404 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    405 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    406 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    407 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    408 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    409 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    410 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    411 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    412 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    413 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    414 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    415 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    416 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    417 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    418 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    419 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    420 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    421 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    422 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    423 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    424 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    425 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    426 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    427 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    428 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    429 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    430 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    431 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    432 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    433 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    434 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    435 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    436 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    437 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    438 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    439 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    440 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    441 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    442 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    443 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    444 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    445 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    446 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    447 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    448 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    449 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    450 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    451 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    452 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    453 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    454 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    455 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    456 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    457 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    458 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    459 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    460 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    461 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    462 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    463 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    464 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    465 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    466 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    467 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    468 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    469 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    470 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    471 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    472 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    473 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    474 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    475 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    476 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    477 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    478 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    479 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    480 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    481 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    482 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    483 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    484 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    485 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    486 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    487 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    488 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    489 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    490 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    491 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    492 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    493 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    494 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    495 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    496 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    497 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    498 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    499 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    500 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    501 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    502 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    503 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    504 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    505 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    506 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    507 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    508 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    509 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    510 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111",
    511 => "00000000000000000000000000000000000000000000000000000000000111111111000000000000000111111111"
  );

  signal ram : ram_type := INIT_BRAM;

  -- Pipelined outputs
  type pipeline_array is array (0 to LATENCY - 1) of std_logic_vector(DATA_WIDTH - 1 downto 0);
  signal pipeline_a : pipeline_array := (others => (others => '1'));
  signal pipeline_b : pipeline_array := (others => (others => '1'));

begin

  process (clk)
    variable addr_a_int, addr_b_int : integer;
  begin
    if rising_edge(clk) then

      -- Convert addresses
      addr_a_int := to_integer(unsigned(addra));
      addr_b_int := to_integer(unsigned(addrb));

      -- Port A: READ_FIRST
      if ena = '1' then
        -- First capture read value
        pipeline_a(0) <= ram(addr_a_int);
        -- Then perform write (doesn't affect current read output)
        if wea = '1' then
          ram(addr_a_int) <= dia;
        end if;
      end if;

      -- Port B: READ_FIRST
      if enb = '1' then
        pipeline_b(0) <= ram(addr_b_int);
        -- Port B write only if not conflicting
        if web = '1' and not (wea = '1' and addr_a_int = addr_b_int) then
          ram(addr_b_int) <= dib;
        end if;
      end if;

      -- Shift pipelines for latency
      for i in 1 to LATENCY - 1 loop
        pipeline_a(i) <= pipeline_a(i - 1);
        pipeline_b(i) <= pipeline_b(i - 1);
      end loop;

    end if;
  end process;

  -- Outputs after constant latency
  doa <= pipeline_a(LATENCY - 1);
  dob <= pipeline_b(LATENCY - 1);

end architecture;
