library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.NUMERIC_STD.all;
  use work.constants_pkg.all;
  use work.bram_init_pkg.all; -- Import constants

entity pipelined_stack_processor is
  port (
    clk : in std_logic;
    rst : in std_logic
  );
end entity;

architecture rtl of pipelined_stack_processor is

  -- BRAM component declaration
  component Flow_mem is
    generic (
      LATENCY : integer
    );
    port (
      clk          : in  std_logic;
      ena, enb     : in  std_logic;
      wea, web     : in  std_logic;
      addra, addrb : in  std_logic_vector(MEM_ADDR_WIDTH - 1 downto 0);
      dia, dib     : in  std_logic_vector(FLOW_MEM_DATA_WIDTH - 1 downto 0);
      doa, dob     : out std_logic_vector(FLOW_MEM_DATA_WIDTH - 1 downto 0)
    );
  end component;

  component Rate_mem is
    generic (
      LATENCY : integer
    );
    port (
      clk          : in  std_logic;
      ena, enb     : in  std_logic;
      wea, web     : in  std_logic;
      addra, addrb : in  std_logic_vector(MEM_ADDR_WIDTH - 1 downto 0);
      dia, dib     : in  std_logic_vector(RATE_MEM_DATA_WIDTH - 1 downto 0);
      doa, dob     : out std_logic_vector(RATE_MEM_DATA_WIDTH - 1 downto 0)
    );
  end component;

  component Calendar is
    port (
      clk            : in  std_logic;
      rst            : in  std_logic;
      insert_enable  : in  std_logic;
      insert_slot    : in  unsigned(CALENDAR_SLOTS_WIDTH - 1 downto 0);
      insert_address : in  std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0);
      current_slot_o : out unsigned(CALENDAR_SLOTS_WIDTH - 1 downto 0);
      head_address_o : out std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0);
      slot_advance_o : out std_logic -- Pulse when moving to the next slot
    );
  end component;

  constant QP_padding : std_logic_vector(QP_WIDTH - FLOW_ADDRESS_WIDTH - 1 downto 0) := (others => '0'); -- Padding for QP

  -- Pipeline registers
  type pipe_stage is record
    valid       : std_logic;
    --qp          : std_logic_vector(QP_WIDTH - 1 downto 0); qp ommitted in the pipeline, current address is used instead
    cur_addr    : std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0);
    next_addr   : std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0);
    max_rate    : unsigned(RATE_BIT_RESOLUTION_WIDTH - 1 downto 0);
    cur_rate    : unsigned(RATE_BIT_RESOLUTION_WIDTH - 1 downto 0);
    seq_nr      : unsigned(SEQ_NR_WIDTH - 1 downto 0);
    active_flag : std_logic;
    --data        : std_logic_vector(DATA_WIDTH - 1 downto 0);
    --processed : std_logic_vector(DATA_WIDTH - 1 downto 0);
  end record;

  type pipe_type is array (0 to PIPELINE_SIZE - 1) of pipe_stage;

  signal pipe_valid : std_logic_vector(PIPELINE_SIZE - 1 downto 0) := (others => '0');
  signal pipe       : pipe_type                                    := (others => (valid => '0', cur_addr => FLOW_NULL_ADDRESS, next_addr => FLOW_NULL_ADDRESS, max_rate => (others => '0'), cur_rate => (others => '0'), seq_nr => (others => '0'), active_flag => '0'));

  -- Internal flow_mem signals
  signal flow_mem_ena   : std_logic                                          := '0';
  signal flow_mem_wea   : std_logic                                          := '0';
  signal flow_mem_addra : std_logic_vector(MEM_ADDR_WIDTH - 1 downto 0)      := MEM_DEFAULT_ADDRESS;
  signal flow_mem_dia   : std_logic_vector(FLOW_MEM_DATA_WIDTH - 1 downto 0) := (others => '0');
  signal flow_mem_doa   : std_logic_vector(FLOW_MEM_DATA_WIDTH - 1 downto 0) := (others => '0');

  signal rate_mem_ena   : std_logic                                          := '0';
  signal rate_mem_wea   : std_logic                                          := '0';
  signal rate_mem_addra : std_logic_vector(MEM_ADDR_WIDTH - 1 downto 0)      := MEM_DEFAULT_ADDRESS;
  signal rate_mem_dia   : std_logic_vector(RATE_MEM_DATA_WIDTH - 1 downto 0) := (others => '0');
  signal rate_mem_doa   : std_logic_vector(RATE_MEM_DATA_WIDTH - 1 downto 0) := (others => '0');

  -- Calendar signals
  signal insert_enable  : std_logic                                         := '0';
  signal insert_slot    : unsigned(CALENDAR_SLOTS_WIDTH - 1 downto 0)       := (others => '0');
  signal insert_address : std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0) := (others => '0');
  signal current_slot_o : unsigned(CALENDAR_SLOTS_WIDTH - 1 downto 0);
  signal head_address_o : std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0);
  signal slot_advance_o : std_logic;
  signal target_slot    : unsigned(CALENDAR_SLOTS_WIDTH - 1 downto 0)       := (others => '0');

begin

  -- Instantiate the BRAM internally
  flow_mem_inst: Flow_mem
    generic map (
      LATENCY => MEM_LATENCY
    )
    port map (
      clk   => clk,
      ena   => flow_mem_ena,
      wea   => flow_mem_wea,
      addra => flow_mem_addra,
      dia   => flow_mem_dia,
      doa   => flow_mem_doa,
      enb   => '0',
      web   => '0',
      addrb => MEM_DEFAULT_ADDRESS,
      dib   => (others => '0'),
      dob   => open
    );

  rate_mem_inst: Rate_mem
    generic map (
      LATENCY => MEM_LATENCY
    )
    port map (
      clk   => clk,
      ena   => rate_mem_ena,
      wea   => rate_mem_wea,
      addra => rate_mem_addra,
      dia   => rate_mem_dia,
      doa   => rate_mem_doa,
      enb   => '0',
      web   => '0',
      addrb => MEM_DEFAULT_ADDRESS,
      dib   => (others => '0'),
      dob   => open
    );

  -- Instantiate Calendar
  calendar_inst: Calendar
    port map (
      clk            => clk,
      rst            => rst,
      insert_enable  => insert_enable,
      insert_slot    => insert_slot,
      insert_address => insert_address,
      current_slot_o => current_slot_o,
      head_address_o => head_address_o,
      slot_advance_o => slot_advance_o
    );

  -- Main pipeline logic
  process (clk)
  begin

    if rising_edge(clk) then

      -- Shift pipeline stages
      for i in PIPELINE_SIZE - 1 downto 1 loop
        pipe(i) <= pipe(i - 1);
        pipe_valid(i) <= pipe_valid(i - 1);
      end loop;

      -- Stage 0: input address or feedback
      if slot_advance_o = '1' then
        if head_address_o /= FLOW_NULL_ADDRESS then
          pipe(0).cur_addr <= head_address_o;
          pipe_valid(0) <= '1';
        end if;
      elsif pipe_valid(MEM_LATENCY + 2) = '1' and pipe(MEM_LATENCY + 2).next_addr /= FLOW_NULL_ADDRESS then
        pipe(0).cur_addr <= pipe(MEM_LATENCY + 2).next_addr;
        pipe_valid(0) <= '1';
      else
        pipe_valid(0) <= '0';
      end if;

      -- Stage 0 issues address to both BRAMs
      if pipe_valid(0) = '1' then
        flow_mem_ena <= '1';
        flow_mem_wea <= '0';
        flow_mem_addra <= std_logic_vector(resize(unsigned(pipe(0).cur_addr(MEM_ADDR_WIDTH - 1 downto 0)), MEM_ADDR_WIDTH));

        rate_mem_ena <= '1';
        rate_mem_wea <= '0';
        rate_mem_addra <= std_logic_vector(resize(unsigned(pipe(0).cur_addr(MEM_ADDR_WIDTH - 1 downto 0)), MEM_ADDR_WIDTH));
      else
        flow_mem_ena <= '0';
        rate_mem_ena <= '0';
      end if;

      -- Stage 3: BRAMs data arrives
      -- The flow_mem data is expected to be in the format:
      -- msb -> lsb
      -- [active_flag, seq_nr, next_addr, cur_addr]
      -- [ 1, SEQ_NR_WIDTH, FLOW_ADDRESS_WIDTH, QP_WIDTH[empty bits: QP_padding, FLOW_ADDRESS_WIDTH]]

      -- The rate_mem data is expected to be in the format:
      -- msb -> lsb
      -- [cur_rate, max_rate]
      -- [RATE_BIT_RESOLUTION_WIDTH, RATE_BIT_RESOLUTION_WIDTH]
      if pipe_valid(MEM_LATENCY + 1) = '1' then
        pipe(MEM_LATENCY + 2).cur_addr <= flow_mem_doa(FLOW_ADDRESS_WIDTH - 1 downto 0);
        pipe(MEM_LATENCY + 2).next_addr <= flow_mem_doa(FLOW_ADDRESS_WIDTH + QP_WIDTH - 1 downto QP_WIDTH);
        pipe(MEM_LATENCY + 2).seq_nr <= unsigned(flow_mem_doa(FLOW_ADDRESS_WIDTH + QP_WIDTH + SEQ_NR_WIDTH - 1 downto FLOW_ADDRESS_WIDTH + QP_WIDTH));
        pipe(MEM_LATENCY + 2).active_flag <= flow_mem_doa(FLOW_ADDRESS_WIDTH + QP_WIDTH + SEQ_NR_WIDTH);

        pipe(MEM_LATENCY + 2).max_rate <= unsigned(rate_mem_doa(RATE_BIT_RESOLUTION_WIDTH - 1 downto 0));
        pipe(MEM_LATENCY + 2).cur_rate <= unsigned(rate_mem_doa(2 * RATE_BIT_RESOLUTION_WIDTH - 1 downto RATE_BIT_RESOLUTION_WIDTH));

      end if;

      -- Stage 4: process 1
      if pipe_valid(MEM_LATENCY + 2) = '1' then
        pipe(MEM_LATENCY + 3).seq_nr <= pipe(MEM_LATENCY + 2).seq_nr + 1;
        target_slot <= (current_slot_o + pipe(MEM_LATENCY + 2).cur_rate) and to_unsigned(CALENDAR_SLOTS - 1, CALENDAR_SLOTS_WIDTH); -- schedule in a circular manner
      end if;

      if pipe_valid(MEM_LATENCY + 3) = '1' then
        insert_enable <= '1';
        insert_slot <= target_slot;
        insert_address <= pipe(MEM_LATENCY + 3).cur_addr;
      else
        insert_enable <= '0';
      end if;

      -- Stage 6: writeback
      if pipe_valid(MEM_LATENCY + 4) = '1' then
        flow_mem_ena <= '1';
        flow_mem_wea <= '1';
        flow_mem_addra <= std_logic_vector(resize(unsigned(pipe(MEM_LATENCY + 4).cur_addr(MEM_ADDR_WIDTH - 1 downto 0)), MEM_ADDR_WIDTH));
        flow_mem_dia <= pipe(MEM_LATENCY + 4).active_flag & std_logic_vector(pipe(MEM_LATENCY + 4).seq_nr) & pipe(MEM_LATENCY + 4).next_addr & QP_padding & pipe(MEM_LATENCY + 4).cur_addr;

        rate_mem_ena <= '1';
        rate_mem_wea <= '1';
        rate_mem_addra <= std_logic_vector(resize(unsigned(pipe(MEM_LATENCY + 4).cur_addr(MEM_ADDR_WIDTH - 1 downto 0)), MEM_ADDR_WIDTH));
        rate_mem_dia <= std_logic_vector(pipe(MEM_LATENCY + 4).cur_rate) & std_logic_vector(pipe(MEM_LATENCY + 4).max_rate);

      else
        flow_mem_wea <= '0';
        rate_mem_wea <= '0';
      end if;

      if rst = '1' then
        pipe_valid <= (others => '0');
        flow_mem_ena <= '0';
        flow_mem_wea <= '0';
        flow_mem_addra <= MEM_DEFAULT_ADDRESS;
        flow_mem_dia <= (others => '0');

        rate_mem_ena <= '0';
        rate_mem_wea <= '0';
        rate_mem_addra <= MEM_DEFAULT_ADDRESS;
        rate_mem_dia <= (others => '0');
      end if;

    end if;
  end process;

end architecture;
