-- RP simulation package
library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use ieee.numeric_std.all;
  use work.constants_pkg.all; -- Import constants

package bram_init_pkg is

  -- Memory
  type rate_mem_type is array (0 to 2 ** 4 - 1) of std_logic_vector(3 - 1 downto 0);
  type RP_mem_type is array (0 to 2 ** 4 - 1) of std_logic_vector(105 - 1 downto 0);

  constant init_rate_mem_16 : rate_mem_type := (
    0  => "111",
    1  => "111",
    2  => "111",
    3  => "111",
    4  => "111",
    5  => "111",
    6  => "111",
    7  => "111",
    8  => "111",
    9  => "110",
    10 => "110",
    11 => "110",
    --11 => "100001", -- Test values for scheduler
    12 => "111",
    13 => "111",
    14 => "111",
    15 => "111"
  );

  constant init_RP_mem_16 : RP_mem_type := (
    0  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    1  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    2  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    3  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    4  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    5  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    6  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    7  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    8  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    9  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    10 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    11 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    12 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    13 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    14 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    15 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111"
  );

end package;
