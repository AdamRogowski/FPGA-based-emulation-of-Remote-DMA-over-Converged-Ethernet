library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use ieee.numeric_std.all;
  use work.constants_pkg.all; -- Import constants

package bram_init_pkg is

  -- Memory
  type flow_mem_type is array (0 to 2 ** 10 - 1) of std_logic_vector(47 - 1 downto 0);
  type rate_mem_type is array (0 to 2 ** 10 - 1) of std_logic_vector(9 - 1 downto 0);
  type calendar_mem_type is array (0 to 2 ** 9 - 1) of std_logic_vector(11 - 1 downto 0);

  -- Flow memory data format
  --|active_flag|seq_nr|next_addr|QP|
  --|    1      |   24  |    11    | 11|
  constant init_flow_mem_1024 : flow_mem_type := (
    0    => "10000000000000000000000001111111111100000000000", -- 1, 0
    1    => "10000000000000000000000000000000001000000000001", -- 2, 1
    2    => "10000000000000000000000000000000001100000000010", -- 3, 2
    3    => "10000000000000000000000000000000010000000000011", -- 4, 3
    4    => "10000000000000000000000000000000010100000000100", -- 5, 4
    5    => "10000000000000000000000000000000011000000000101", -- 6, 5
    6    => "10000000000000000000000000000000011100000000110", -- 7, 6
    7    => "10000000000000000000000000000000100000000000111", -- 8, 7
    8    => "10000000000000000000000000000000100100000001000", -- 9, 8
    9    => "10000000000000000000000000000000101000000001001", -- 10, 9
    10   => "10000000000000000000000000000000101100000001010", -- 11, 10
    11   => "10000000000000000000000000000000110000000001011", -- 12, 11
    12   => "10000000000000000000000000000000110100000001100", -- 13, 12
    13   => "10000000000000000000000000000000111000000001101", -- 14, 13
    14   => "10000000000000000000000000000000111100000001110", -- 15, 14
    15   => "10000000000000000000000000000001000000000001111", -- 16, 15
    16   => "10000000000000000000000000000001000100000010000", -- 17, 16
    17   => "10000000000000000000000000000001001000000010001", -- 18, 17
    18   => "10000000000000000000000000000001001100000010010", -- 19, 18
    19   => "10000000000000000000000000000001010000000010011", -- 20, 19
    20   => "10000000000000000000000000000001010100000010100", -- 21, 20
    21   => "10000000000000000000000000000001011000000010101", -- 22, 21
    22   => "10000000000000000000000000000001011100000010110", -- 23, 22
    23   => "10000000000000000000000000000001100000000010111", -- 24, 23
    24   => "10000000000000000000000000000001100100000011000", -- 25, 24
    25   => "10000000000000000000000000000001101000000011001", -- 26, 25
    26   => "10000000000000000000000000000001101100000011010", -- 27, 26
    27   => "10000000000000000000000000000001110000000011011", -- 28, 27
    28   => "10000000000000000000000000000001110100000011100", -- 29, 28
    29   => "10000000000000000000000000000001111000000011101", -- 30, 29
    30   => "10000000000000000000000000000001111100000011110", -- 31, 30
    31   => "10000000000000000000000000000010000000000011111", -- 32, 31
    32   => "10000000000000000000000000000010000100000100000", -- 33, 32
    33   => "10000000000000000000000000000010001000000100001", -- 34, 33
    34   => "10000000000000000000000000000010001100000100010", -- 35, 34
    35   => "10000000000000000000000000000010010000000100011", -- 36, 35
    36   => "10000000000000000000000000000010010100000100100", -- 37, 36
    37   => "10000000000000000000000000000010011000000100101", -- 38, 37
    38   => "10000000000000000000000000000010011100000100110", -- 39, 38
    39   => "10000000000000000000000000000010100000000100111", -- 40, 39
    40   => "10000000000000000000000000000010100100000101000", -- 41, 40
    41   => "10000000000000000000000000000010101000000101001", -- 42, 41
    42   => "10000000000000000000000000000010101100000101010", -- 43, 42
    43   => "10000000000000000000000000000010110000000101011", -- 44, 43
    44   => "10000000000000000000000000000010110100000101100", -- 45, 44
    45   => "10000000000000000000000000000010111000000101101", -- 46, 45
    46   => "10000000000000000000000000000010111100000101110", -- 47, 46
    47   => "10000000000000000000000000000011000000000101111", -- 48, 47
    48   => "10000000000000000000000000000011000100000110000", -- 49, 48
    49   => "10000000000000000000000000000011001000000110001", -- 50, 49
    50   => "10000000000000000000000000000011001100000110010", -- 51, 50
    51   => "10000000000000000000000000000011010000000110011", -- 52, 51
    52   => "10000000000000000000000000000011010100000110100", -- 53, 52
    53   => "10000000000000000000000000000011011000000110101", -- 54, 53
    54   => "10000000000000000000000000000011011100000110110", -- 55, 54
    55   => "10000000000000000000000000000011100000000110111", -- 56, 55
    56   => "10000000000000000000000000000011100100000111000", -- 57, 56
    57   => "10000000000000000000000000000011101000000111001", -- 58, 57
    58   => "10000000000000000000000000000011101100000111010", -- 59, 58
    59   => "10000000000000000000000000000011110000000111011", -- 60, 59
    60   => "10000000000000000000000000000011110100000111100", -- 61, 60
    61   => "10000000000000000000000000000011111000000111101", -- 62, 61
    62   => "10000000000000000000000000000011111100000111110", -- 63, 62
    63   => "10000000000000000000000000000100000000000111111", -- 64, 63
    64   => "10000000000000000000000000000100000100001000000", -- 65, 64
    65   => "10000000000000000000000000000100001000001000001", -- 66, 65
    66   => "10000000000000000000000000000100001100001000010", -- 67, 66
    67   => "10000000000000000000000000000100010000001000011", -- 68, 67
    68   => "10000000000000000000000000000100010100001000100", -- 69, 68
    69   => "10000000000000000000000000000100011000001000101", -- 70, 69
    70   => "10000000000000000000000000000100011100001000110", -- 71, 70
    71   => "10000000000000000000000000000100100000001000111", -- 72, 71
    72   => "10000000000000000000000000000100100100001001000", -- 73, 72
    73   => "10000000000000000000000000000100101000001001001", -- 74, 73
    74   => "10000000000000000000000000000100101100001001010", -- 75, 74
    75   => "10000000000000000000000000000100110000001001011", -- 76, 75
    76   => "10000000000000000000000000000100110100001001100", -- 77, 76
    77   => "10000000000000000000000000000100111000001001101", -- 78, 77
    78   => "10000000000000000000000000000100111100001001110", -- 79, 78
    79   => "10000000000000000000000000000101000000001001111", -- 80, 79
    80   => "10000000000000000000000000000101000100001010000", -- 81, 80
    81   => "10000000000000000000000000000101001000001010001", -- 82, 81
    82   => "10000000000000000000000000000101001100001010010", -- 83, 82
    83   => "10000000000000000000000000000101010000001010011", -- 84, 83
    84   => "10000000000000000000000000000101010100001010100", -- 85, 84
    85   => "10000000000000000000000000000101011000001010101", -- 86, 85
    86   => "10000000000000000000000000000101011100001010110", -- 87, 86
    87   => "10000000000000000000000000000101100000001010111", -- 88, 87
    88   => "10000000000000000000000000000101100100001011000", -- 89, 88
    89   => "10000000000000000000000000000101101000001011001", -- 90, 89
    90   => "10000000000000000000000000000101101100001011010", -- 91, 90
    91   => "10000000000000000000000000000101110000001011011", -- 92, 91
    92   => "10000000000000000000000000000101110100001011100", -- 93, 92
    93   => "10000000000000000000000000000101111000001011101", -- 94, 93
    94   => "10000000000000000000000000000101111100001011110", -- 95, 94
    95   => "10000000000000000000000000000110000000001011111", -- 96, 95
    96   => "10000000000000000000000000000110000100001100000", -- 97, 96
    97   => "10000000000000000000000000000110001000001100001", -- 98, 97
    98   => "10000000000000000000000000000110001100001100010", -- 99, 98
    99   => "10000000000000000000000000000110010000001100011", -- 100, 99
    100  => "10000000000000000000000000000110010100001100100", -- 101, 100
    101  => "10000000000000000000000000000110011000001100101", -- 102, 101
    102  => "10000000000000000000000000000110011100001100110", -- 103, 102
    103  => "10000000000000000000000000000110100000001100111", -- 104, 103
    104  => "10000000000000000000000000000110100100001101000", -- 105, 104
    105  => "10000000000000000000000000000110101000001101001", -- 106, 105
    106  => "10000000000000000000000000000110101100001101010", -- 107, 106
    107  => "10000000000000000000000000000110110000001101011", -- 108, 107
    108  => "10000000000000000000000000000110110100001101100", -- 109, 108
    109  => "10000000000000000000000000000110111000001101101", -- 110, 109
    110  => "10000000000000000000000000000110111100001101110", -- 111, 110
    111  => "10000000000000000000000000000111000000001101111", -- 112, 111
    112  => "10000000000000000000000000000111000100001110000", -- 113, 112
    113  => "10000000000000000000000000000111001000001110001", -- 114, 113
    114  => "10000000000000000000000000000111001100001110010", -- 115, 114
    115  => "10000000000000000000000000000111010000001110011", -- 116, 115
    116  => "10000000000000000000000000000111010100001110100", -- 117, 116
    117  => "10000000000000000000000000000111011000001110101", -- 118, 117
    118  => "10000000000000000000000000000111011100001110110", -- 119, 118
    119  => "10000000000000000000000000000111100000001110111", -- 120, 119
    120  => "10000000000000000000000000000111100100001111000", -- 121, 120
    121  => "10000000000000000000000000000111101000001111001", -- 122, 121
    122  => "10000000000000000000000000000111101100001111010", -- 123, 122
    123  => "10000000000000000000000000000111110000001111011", -- 124, 123
    124  => "10000000000000000000000000000111110100001111100", -- 125, 124
    125  => "10000000000000000000000000000111111000001111101", -- 126, 125
    126  => "10000000000000000000000000000111111100001111110", -- 127, 126
    127  => "10000000000000000000000000001000000000001111111", -- 128, 127
    128  => "10000000000000000000000000001000000100010000000", -- 129, 128
    129  => "10000000000000000000000000001000001000010000001", -- 130, 129
    130  => "10000000000000000000000000001000001100010000010", -- 131, 130
    131  => "10000000000000000000000000001000010000010000011", -- 132, 131
    132  => "10000000000000000000000000001000010100010000100", -- 133, 132
    133  => "10000000000000000000000000001000011000010000101", -- 134, 133
    134  => "10000000000000000000000000001000011100010000110", -- 135, 134
    135  => "10000000000000000000000000001000100000010000111", -- 136, 135
    136  => "10000000000000000000000000001000100100010001000", -- 137, 136
    137  => "10000000000000000000000000001000101000010001001", -- 138, 137
    138  => "10000000000000000000000000001000101100010001010", -- 139, 138
    139  => "10000000000000000000000000001000110000010001011", -- 140, 139
    140  => "10000000000000000000000000001000110100010001100", -- 141, 140
    141  => "10000000000000000000000000001000111000010001101", -- 142, 141
    142  => "10000000000000000000000000001000111100010001110", -- 143, 142
    143  => "10000000000000000000000000001001000000010001111", -- 144, 143
    144  => "10000000000000000000000000001001000100010010000", -- 145, 144
    145  => "10000000000000000000000000001001001000010010001", -- 146, 145
    146  => "10000000000000000000000000001001001100010010010", -- 147, 146
    147  => "10000000000000000000000000001001010000010010011", -- 148, 147
    148  => "10000000000000000000000000001001010100010010100", -- 149, 148
    149  => "10000000000000000000000000001001011000010010101", -- 150, 149
    150  => "10000000000000000000000000001001011100010010110", -- 151, 150
    151  => "10000000000000000000000000001001100000010010111", -- 152, 151
    152  => "10000000000000000000000000001001100100010011000", -- 153, 152
    153  => "10000000000000000000000000001001101000010011001", -- 154, 153
    154  => "10000000000000000000000000001001101100010011010", -- 155, 154
    155  => "10000000000000000000000000001001110000010011011", -- 156, 155
    156  => "10000000000000000000000000001001110100010011100", -- 157, 156
    157  => "10000000000000000000000000001001111000010011101", -- 158, 157
    158  => "10000000000000000000000000001001111100010011110", -- 159, 158
    159  => "10000000000000000000000000001010000000010011111", -- 160, 159
    160  => "10000000000000000000000000001010000100010100000", -- 161, 160
    161  => "10000000000000000000000000001010001000010100001", -- 162, 161
    162  => "10000000000000000000000000001010001100010100010", -- 163, 162
    163  => "10000000000000000000000000001010010000010100011", -- 164, 163
    164  => "10000000000000000000000000001010010100010100100", -- 165, 164
    165  => "10000000000000000000000000001010011000010100101", -- 166, 165
    166  => "10000000000000000000000000001010011100010100110", -- 167, 166
    167  => "10000000000000000000000000001010100000010100111", -- 168, 167
    168  => "10000000000000000000000000001010100100010101000", -- 169, 168
    169  => "10000000000000000000000000001010101000010101001", -- 170, 169
    170  => "10000000000000000000000000001010101100010101010", -- 171, 170
    171  => "10000000000000000000000000001010110000010101011", -- 172, 171
    172  => "10000000000000000000000000001010110100010101100", -- 173, 172
    173  => "10000000000000000000000000001010111000010101101", -- 174, 173
    174  => "10000000000000000000000000001010111100010101110", -- 175, 174
    175  => "10000000000000000000000000001011000000010101111", -- 176, 175
    176  => "10000000000000000000000000001011000100010110000", -- 177, 176
    177  => "10000000000000000000000000001011001000010110001", -- 178, 177
    178  => "10000000000000000000000000001011001100010110010", -- 179, 178
    179  => "10000000000000000000000000001011010000010110011", -- 180, 179
    180  => "10000000000000000000000000001011010100010110100", -- 181, 180
    181  => "10000000000000000000000000001011011000010110101", -- 182, 181
    182  => "10000000000000000000000000001011011100010110110", -- 183, 182
    183  => "10000000000000000000000000001011100000010110111", -- 184, 183
    184  => "10000000000000000000000000001011100100010111000", -- 185, 184
    185  => "10000000000000000000000000001011101000010111001", -- 186, 185
    186  => "10000000000000000000000000001011101100010111010", -- 187, 186
    187  => "10000000000000000000000000001011110000010111011", -- 188, 187
    188  => "10000000000000000000000000001011110100010111100", -- 189, 188
    189  => "10000000000000000000000000001011111000010111101", -- 190, 189
    190  => "10000000000000000000000000001011111100010111110", -- 191, 190
    191  => "10000000000000000000000000001100000000010111111", -- 192, 191
    192  => "10000000000000000000000000001100000100011000000", -- 193, 192
    193  => "10000000000000000000000000001100001000011000001", -- 194, 193
    194  => "10000000000000000000000000001100001100011000010", -- 195, 194
    195  => "10000000000000000000000000001100010000011000011", -- 196, 195
    196  => "10000000000000000000000000001100010100011000100", -- 197, 196
    197  => "10000000000000000000000000001100011000011000101", -- 198, 197
    198  => "10000000000000000000000000001100011100011000110", -- 199, 198
    199  => "10000000000000000000000000001100100000011000111", -- 200, 199
    200  => "10000000000000000000000000001100100100011001000", -- 201, 200
    201  => "10000000000000000000000000001100101000011001001", -- 202, 201
    202  => "10000000000000000000000000001100101100011001010", -- 203, 202
    203  => "10000000000000000000000000001100110000011001011", -- 204, 203
    204  => "10000000000000000000000000001100110100011001100", -- 205, 204
    205  => "10000000000000000000000000001100111000011001101", -- 206, 205
    206  => "10000000000000000000000000001100111100011001110", -- 207, 206
    207  => "10000000000000000000000000001101000000011001111", -- 208, 207
    208  => "10000000000000000000000000001101000100011010000", -- 209, 208
    209  => "10000000000000000000000000001101001000011010001", -- 210, 209
    210  => "10000000000000000000000000001101001100011010010", -- 211, 210
    211  => "10000000000000000000000000001101010000011010011", -- 212, 211
    212  => "10000000000000000000000000001101010100011010100", -- 213, 212
    213  => "10000000000000000000000000001101011000011010101", -- 214, 213
    214  => "10000000000000000000000000001101011100011010110", -- 215, 214
    215  => "10000000000000000000000000001101100000011010111", -- 216, 215
    216  => "10000000000000000000000000001101100100011011000", -- 217, 216
    217  => "10000000000000000000000000001101101000011011001", -- 218, 217
    218  => "10000000000000000000000000001101101100011011010", -- 219, 218
    219  => "10000000000000000000000000001101110000011011011", -- 220, 219
    220  => "10000000000000000000000000001101110100011011100", -- 221, 220
    221  => "10000000000000000000000000001101111000011011101", -- 222, 221
    222  => "10000000000000000000000000001101111100011011110", -- 223, 222
    223  => "10000000000000000000000000001110000000011011111", -- 224, 223
    224  => "10000000000000000000000000001110000100011100000", -- 225, 224
    225  => "10000000000000000000000000001110001000011100001", -- 226, 225
    226  => "10000000000000000000000000001110001100011100010", -- 227, 226
    227  => "10000000000000000000000000001110010000011100011", -- 228, 227
    228  => "10000000000000000000000000001110010100011100100", -- 229, 228
    229  => "10000000000000000000000000001110011000011100101", -- 230, 229
    230  => "10000000000000000000000000001110011100011100110", -- 231, 230
    231  => "10000000000000000000000000001110100000011100111", -- 232, 231
    232  => "10000000000000000000000000001110100100011101000", -- 233, 232
    233  => "10000000000000000000000000001110101000011101001", -- 234, 233
    234  => "10000000000000000000000000001110101100011101010", -- 235, 234
    235  => "10000000000000000000000000001110110000011101011", -- 236, 235
    236  => "10000000000000000000000000001110110100011101100", -- 237, 236
    237  => "10000000000000000000000000001110111000011101101", -- 238, 237
    238  => "10000000000000000000000000001110111100011101110", -- 239, 238
    239  => "10000000000000000000000000001111000000011101111", -- 240, 239
    240  => "10000000000000000000000000001111000100011110000", -- 241, 240
    241  => "10000000000000000000000000001111001000011110001", -- 242, 241
    242  => "10000000000000000000000000001111001100011110010", -- 243, 242
    243  => "10000000000000000000000000001111010000011110011", -- 244, 243
    244  => "10000000000000000000000000001111010100011110100", -- 245, 244
    245  => "10000000000000000000000000001111011000011110101", -- 246, 245
    246  => "10000000000000000000000000001111011100011110110", -- 247, 246
    247  => "10000000000000000000000000001111100000011110111", -- 248, 247
    248  => "10000000000000000000000000001111100100011111000", -- 249, 248
    249  => "10000000000000000000000000001111101000011111001", -- 250, 249
    250  => "10000000000000000000000000001111101100011111010", -- 251, 250
    251  => "10000000000000000000000000001111110000011111011", -- 252, 251
    252  => "10000000000000000000000000001111110100011111100", -- 253, 252
    253  => "10000000000000000000000000001111111000011111101", -- 254, 253
    254  => "10000000000000000000000000001111111100011111110", -- 255, 254
    255  => "10000000000000000000000000010000000000011111111", -- 256, 255
    256  => "10000000000000000000000000010000000100100000000", -- 257, 256
    257  => "10000000000000000000000000010000001000100000001", -- 258, 257
    258  => "10000000000000000000000000010000001100100000010", -- 259, 258
    259  => "10000000000000000000000000010000010000100000011", -- 260, 259
    260  => "10000000000000000000000000010000010100100000100", -- 261, 260
    261  => "10000000000000000000000000010000011000100000101", -- 262, 261
    262  => "10000000000000000000000000010000011100100000110", -- 263, 262
    263  => "10000000000000000000000000010000100000100000111", -- 264, 263
    264  => "10000000000000000000000000010000100100100001000", -- 265, 264
    265  => "10000000000000000000000000010000101000100001001", -- 266, 265
    266  => "10000000000000000000000000010000101100100001010", -- 267, 266
    267  => "10000000000000000000000000010000110000100001011", -- 268, 267
    268  => "10000000000000000000000000010000110100100001100", -- 269, 268
    269  => "10000000000000000000000000010000111000100001101", -- 270, 269
    270  => "10000000000000000000000000010000111100100001110", -- 271, 270
    271  => "10000000000000000000000000010001000000100001111", -- 272, 271
    272  => "10000000000000000000000000010001000100100010000", -- 273, 272
    273  => "10000000000000000000000000010001001000100010001", -- 274, 273
    274  => "10000000000000000000000000010001001100100010010", -- 275, 274
    275  => "10000000000000000000000000010001010000100010011", -- 276, 275
    276  => "10000000000000000000000000010001010100100010100", -- 277, 276
    277  => "10000000000000000000000000010001011000100010101", -- 278, 277
    278  => "10000000000000000000000000010001011100100010110", -- 279, 278
    279  => "10000000000000000000000000010001100000100010111", -- 280, 279
    280  => "10000000000000000000000000010001100100100011000", -- 281, 280
    281  => "10000000000000000000000000010001101000100011001", -- 282, 281
    282  => "10000000000000000000000000010001101100100011010", -- 283, 282
    283  => "10000000000000000000000000010001110000100011011", -- 284, 283
    284  => "10000000000000000000000000010001110100100011100", -- 285, 284
    285  => "10000000000000000000000000010001111000100011101", -- 286, 285
    286  => "10000000000000000000000000010001111100100011110", -- 287, 286
    287  => "10000000000000000000000000010010000000100011111", -- 288, 287
    288  => "10000000000000000000000000010010000100100100000", -- 289, 288
    289  => "10000000000000000000000000010010001000100100001", -- 290, 289
    290  => "10000000000000000000000000010010001100100100010", -- 291, 290
    291  => "10000000000000000000000000010010010000100100011", -- 292, 291
    292  => "10000000000000000000000000010010010100100100100", -- 293, 292
    293  => "10000000000000000000000000010010011000100100101", -- 294, 293
    294  => "10000000000000000000000000010010011100100100110", -- 295, 294
    295  => "10000000000000000000000000010010100000100100111", -- 296, 295
    296  => "10000000000000000000000000010010100100100101000", -- 297, 296
    297  => "10000000000000000000000000010010101000100101001", -- 298, 297
    298  => "10000000000000000000000000010010101100100101010", -- 299, 298
    299  => "10000000000000000000000000010010110000100101011", -- 300, 299
    300  => "10000000000000000000000000010010110100100101100", -- 301, 300
    301  => "10000000000000000000000000010010111000100101101", -- 302, 301
    302  => "10000000000000000000000000010010111100100101110", -- 303, 302
    303  => "10000000000000000000000000010011000000100101111", -- 304, 303
    304  => "10000000000000000000000000010011000100100110000", -- 305, 304
    305  => "10000000000000000000000000010011001000100110001", -- 306, 305
    306  => "10000000000000000000000000010011001100100110010", -- 307, 306
    307  => "10000000000000000000000000010011010000100110011", -- 308, 307
    308  => "10000000000000000000000000010011010100100110100", -- 309, 308
    309  => "10000000000000000000000000010011011000100110101", -- 310, 309
    310  => "10000000000000000000000000010011011100100110110", -- 311, 310
    311  => "10000000000000000000000000010011100000100110111", -- 312, 311
    312  => "10000000000000000000000000010011100100100111000", -- 313, 312
    313  => "10000000000000000000000000010011101000100111001", -- 314, 313
    314  => "10000000000000000000000000010011101100100111010", -- 315, 314
    315  => "10000000000000000000000000010011110000100111011", -- 316, 315
    316  => "10000000000000000000000000010011110100100111100", -- 317, 316
    317  => "10000000000000000000000000010011111000100111101", -- 318, 317
    318  => "10000000000000000000000000010011111100100111110", -- 319, 318
    319  => "10000000000000000000000000010100000000100111111", -- 320, 319
    320  => "10000000000000000000000000010100000100101000000", -- 321, 320
    321  => "10000000000000000000000000010100001000101000001", -- 322, 321
    322  => "10000000000000000000000000010100001100101000010", -- 323, 322
    323  => "10000000000000000000000000010100010000101000011", -- 324, 323
    324  => "10000000000000000000000000010100010100101000100", -- 325, 324
    325  => "10000000000000000000000000010100011000101000101", -- 326, 325
    326  => "10000000000000000000000000010100011100101000110", -- 327, 326
    327  => "10000000000000000000000000010100100000101000111", -- 328, 327
    328  => "10000000000000000000000000010100100100101001000", -- 329, 328
    329  => "10000000000000000000000000010100101000101001001", -- 330, 329
    330  => "10000000000000000000000000010100101100101001010", -- 331, 330
    331  => "10000000000000000000000000010100110000101001011", -- 332, 331
    332  => "10000000000000000000000000010100110100101001100", -- 333, 332
    333  => "10000000000000000000000000010100111000101001101", -- 334, 333
    334  => "10000000000000000000000000010100111100101001110", -- 335, 334
    335  => "10000000000000000000000000010101000000101001111", -- 336, 335
    336  => "10000000000000000000000000010101000100101010000", -- 337, 336
    337  => "10000000000000000000000000010101001000101010001", -- 338, 337
    338  => "10000000000000000000000000010101001100101010010", -- 339, 338
    339  => "10000000000000000000000000010101010000101010011", -- 340, 339
    340  => "10000000000000000000000000010101010100101010100", -- 341, 340
    341  => "10000000000000000000000000010101011000101010101", -- 342, 341
    342  => "10000000000000000000000000010101011100101010110", -- 343, 342
    343  => "10000000000000000000000000010101100000101010111", -- 344, 343
    344  => "10000000000000000000000000010101100100101011000", -- 345, 344
    345  => "10000000000000000000000000010101101000101011001", -- 346, 345
    346  => "10000000000000000000000000010101101100101011010", -- 347, 346
    347  => "10000000000000000000000000010101110000101011011", -- 348, 347
    348  => "10000000000000000000000000010101110100101011100", -- 349, 348
    349  => "10000000000000000000000000010101111000101011101", -- 350, 349
    350  => "10000000000000000000000000010101111100101011110", -- 351, 350
    351  => "10000000000000000000000000010110000000101011111", -- 352, 351
    352  => "10000000000000000000000000010110000100101100000", -- 353, 352
    353  => "10000000000000000000000000010110001000101100001", -- 354, 353
    354  => "10000000000000000000000000010110001100101100010", -- 355, 354
    355  => "10000000000000000000000000010110010000101100011", -- 356, 355
    356  => "10000000000000000000000000010110010100101100100", -- 357, 356
    357  => "10000000000000000000000000010110011000101100101", -- 358, 357
    358  => "10000000000000000000000000010110011100101100110", -- 359, 358
    359  => "10000000000000000000000000010110100000101100111", -- 360, 359
    360  => "10000000000000000000000000010110100100101101000", -- 361, 360
    361  => "10000000000000000000000000010110101000101101001", -- 362, 361
    362  => "10000000000000000000000000010110101100101101010", -- 363, 362
    363  => "10000000000000000000000000010110110000101101011", -- 364, 363
    364  => "10000000000000000000000000010110110100101101100", -- 365, 364
    365  => "10000000000000000000000000010110111000101101101", -- 366, 365
    366  => "10000000000000000000000000010110111100101101110", -- 367, 366
    367  => "10000000000000000000000000010111000000101101111", -- 368, 367
    368  => "10000000000000000000000000010111000100101110000", -- 369, 368
    369  => "10000000000000000000000000010111001000101110001", -- 370, 369
    370  => "10000000000000000000000000010111001100101110010", -- 371, 370
    371  => "10000000000000000000000000010111010000101110011", -- 372, 371
    372  => "10000000000000000000000000010111010100101110100", -- 373, 372
    373  => "10000000000000000000000000010111011000101110101", -- 374, 373
    374  => "10000000000000000000000000010111011100101110110", -- 375, 374
    375  => "10000000000000000000000000010111100000101110111", -- 376, 375
    376  => "10000000000000000000000000010111100100101111000", -- 377, 376
    377  => "10000000000000000000000000010111101000101111001", -- 378, 377
    378  => "10000000000000000000000000010111101100101111010", -- 379, 378
    379  => "10000000000000000000000000010111110000101111011", -- 380, 379
    380  => "10000000000000000000000000010111110100101111100", -- 381, 380
    381  => "10000000000000000000000000010111111000101111101", -- 382, 381
    382  => "10000000000000000000000000010111111100101111110", -- 383, 382
    383  => "10000000000000000000000000011000000000101111111", -- 384, 383
    384  => "10000000000000000000000000011000000100110000000", -- 385, 384
    385  => "10000000000000000000000000011000001000110000001", -- 386, 385
    386  => "10000000000000000000000000011000001100110000010", -- 387, 386
    387  => "10000000000000000000000000011000010000110000011", -- 388, 387
    388  => "10000000000000000000000000011000010100110000100", -- 389, 388
    389  => "10000000000000000000000000011000011000110000101", -- 390, 389
    390  => "10000000000000000000000000011000011100110000110", -- 391, 390
    391  => "10000000000000000000000000011000100000110000111", -- 392, 391
    392  => "10000000000000000000000000011000100100110001000", -- 393, 392
    393  => "10000000000000000000000000011000101000110001001", -- 394, 393
    394  => "10000000000000000000000000011000101100110001010", -- 395, 394
    395  => "10000000000000000000000000011000110000110001011", -- 396, 395
    396  => "10000000000000000000000000011000110100110001100", -- 397, 396
    397  => "10000000000000000000000000011000111000110001101", -- 398, 397
    398  => "10000000000000000000000000011000111100110001110", -- 399, 398
    399  => "10000000000000000000000000011001000000110001111", -- 400, 399
    400  => "10000000000000000000000000011001000100110010000", -- 401, 400
    401  => "10000000000000000000000000011001001000110010001", -- 402, 401
    402  => "10000000000000000000000000011001001100110010010", -- 403, 402
    403  => "10000000000000000000000000011001010000110010011", -- 404, 403
    404  => "10000000000000000000000000011001010100110010100", -- 405, 404
    405  => "10000000000000000000000000011001011000110010101", -- 406, 405
    406  => "10000000000000000000000000011001011100110010110", -- 407, 406
    407  => "10000000000000000000000000011001100000110010111", -- 408, 407
    408  => "10000000000000000000000000011001100100110011000", -- 409, 408
    409  => "10000000000000000000000000011001101000110011001", -- 410, 409
    410  => "10000000000000000000000000011001101100110011010", -- 411, 410
    411  => "10000000000000000000000000011001110000110011011", -- 412, 411
    412  => "10000000000000000000000000011001110100110011100", -- 413, 412
    413  => "10000000000000000000000000011001111000110011101", -- 414, 413
    414  => "10000000000000000000000000011001111100110011110", -- 415, 414
    415  => "10000000000000000000000000011010000000110011111", -- 416, 415
    416  => "10000000000000000000000000011010000100110100000", -- 417, 416
    417  => "10000000000000000000000000011010001000110100001", -- 418, 417
    418  => "10000000000000000000000000011010001100110100010", -- 419, 418
    419  => "10000000000000000000000000011010010000110100011", -- 420, 419
    420  => "10000000000000000000000000011010010100110100100", -- 421, 420
    421  => "10000000000000000000000000011010011000110100101", -- 422, 421
    422  => "10000000000000000000000000011010011100110100110", -- 423, 422
    423  => "10000000000000000000000000011010100000110100111", -- 424, 423
    424  => "10000000000000000000000000011010100100110101000", -- 425, 424
    425  => "10000000000000000000000000011010101000110101001", -- 426, 425
    426  => "10000000000000000000000000011010101100110101010", -- 427, 426
    427  => "10000000000000000000000000011010110000110101011", -- 428, 427
    428  => "10000000000000000000000000011010110100110101100", -- 429, 428
    429  => "10000000000000000000000000011010111000110101101", -- 430, 429
    430  => "10000000000000000000000000011010111100110101110", -- 431, 430
    431  => "10000000000000000000000000011011000000110101111", -- 432, 431
    432  => "10000000000000000000000000011011000100110110000", -- 433, 432
    433  => "10000000000000000000000000011011001000110110001", -- 434, 433
    434  => "10000000000000000000000000011011001100110110010", -- 435, 434
    435  => "10000000000000000000000000011011010000110110011", -- 436, 435
    436  => "10000000000000000000000000011011010100110110100", -- 437, 436
    437  => "10000000000000000000000000011011011000110110101", -- 438, 437
    438  => "10000000000000000000000000011011011100110110110", -- 439, 438
    439  => "10000000000000000000000000011011100000110110111", -- 440, 439
    440  => "10000000000000000000000000011011100100110111000", -- 441, 440
    441  => "10000000000000000000000000011011101000110111001", -- 442, 441
    442  => "10000000000000000000000000011011101100110111010", -- 443, 442
    443  => "10000000000000000000000000011011110000110111011", -- 444, 443
    444  => "10000000000000000000000000011011110100110111100", -- 445, 444
    445  => "10000000000000000000000000011011111000110111101", -- 446, 445
    446  => "10000000000000000000000000011011111100110111110", -- 447, 446
    447  => "10000000000000000000000000011100000000110111111", -- 448, 447
    448  => "10000000000000000000000000011100000100111000000", -- 449, 448
    449  => "10000000000000000000000000011100001000111000001", -- 450, 449
    450  => "10000000000000000000000000011100001100111000010", -- 451, 450
    451  => "10000000000000000000000000011100010000111000011", -- 452, 451
    452  => "10000000000000000000000000011100010100111000100", -- 453, 452
    453  => "10000000000000000000000000011100011000111000101", -- 454, 453
    454  => "10000000000000000000000000011100011100111000110", -- 455, 454
    455  => "10000000000000000000000000011100100000111000111", -- 456, 455
    456  => "10000000000000000000000000011100100100111001000", -- 457, 456
    457  => "10000000000000000000000000011100101000111001001", -- 458, 457
    458  => "10000000000000000000000000011100101100111001010", -- 459, 458
    459  => "10000000000000000000000000011100110000111001011", -- 460, 459
    460  => "10000000000000000000000000011100110100111001100", -- 461, 460
    461  => "10000000000000000000000000011100111000111001101", -- 462, 461
    462  => "10000000000000000000000000011100111100111001110", -- 463, 462
    463  => "10000000000000000000000000011101000000111001111", -- 464, 463
    464  => "10000000000000000000000000011101000100111010000", -- 465, 464
    465  => "10000000000000000000000000011101001000111010001", -- 466, 465
    466  => "10000000000000000000000000011101001100111010010", -- 467, 466
    467  => "10000000000000000000000000011101010000111010011", -- 468, 467
    468  => "10000000000000000000000000011101010100111010100", -- 469, 468
    469  => "10000000000000000000000000011101011000111010101", -- 470, 469
    470  => "10000000000000000000000000011101011100111010110", -- 471, 470
    471  => "10000000000000000000000000011101100000111010111", -- 472, 471
    472  => "10000000000000000000000000011101100100111011000", -- 473, 472
    473  => "10000000000000000000000000011101101000111011001", -- 474, 473
    474  => "10000000000000000000000000011101101100111011010", -- 475, 474
    475  => "10000000000000000000000000011101110000111011011", -- 476, 475
    476  => "10000000000000000000000000011101110100111011100", -- 477, 476
    477  => "10000000000000000000000000011101111000111011101", -- 478, 477
    478  => "10000000000000000000000000011101111100111011110", -- 479, 478
    479  => "10000000000000000000000000011110000000111011111", -- 480, 479
    480  => "10000000000000000000000000011110000100111100000", -- 481, 480
    481  => "10000000000000000000000000011110001000111100001", -- 482, 481
    482  => "10000000000000000000000000011110001100111100010", -- 483, 482
    483  => "10000000000000000000000000011110010000111100011", -- 484, 483
    484  => "10000000000000000000000000011110010100111100100", -- 485, 484
    485  => "10000000000000000000000000011110011000111100101", -- 486, 485
    486  => "10000000000000000000000000011110011100111100110", -- 487, 486
    487  => "10000000000000000000000000011110100000111100111", -- 488, 487
    488  => "10000000000000000000000000011110100100111101000", -- 489, 488
    489  => "10000000000000000000000000011110101000111101001", -- 490, 489
    490  => "10000000000000000000000000011110101100111101010", -- 491, 490
    491  => "10000000000000000000000000011110110000111101011", -- 492, 491
    492  => "10000000000000000000000000011110110100111101100", -- 493, 492
    493  => "10000000000000000000000000011110111000111101101", -- 494, 493
    494  => "10000000000000000000000000011110111100111101110", -- 495, 494
    495  => "10000000000000000000000000011111000000111101111", -- 496, 495
    496  => "10000000000000000000000000011111000100111110000", -- 497, 496
    497  => "10000000000000000000000000011111001000111110001", -- 498, 497
    498  => "10000000000000000000000000011111001100111110010", -- 499, 498
    499  => "10000000000000000000000000011111010000111110011", -- 500, 499
    500  => "10000000000000000000000000011111010100111110100", -- 501, 500
    501  => "10000000000000000000000000011111011000111110101", -- 502, 501
    502  => "10000000000000000000000000011111011100111110110", -- 503, 502
    503  => "10000000000000000000000000011111100000111110111", -- 504, 503
    504  => "10000000000000000000000000011111100100111111000", -- 505, 504
    505  => "10000000000000000000000000011111101000111111001", -- 506, 505
    506  => "10000000000000000000000000011111101100111111010", -- 507, 506
    507  => "10000000000000000000000000011111110000111111011", -- 508, 507
    508  => "10000000000000000000000000011111110100111111100", -- 509, 508
    509  => "10000000000000000000000000011111111000111111101", -- 510, 509
    510  => "10000000000000000000000000011111111100111111110", -- 511, 510
    511  => "10000000000000000000000000100000000000111111111", -- 512, 511
    512  => "10000000000000000000000000100000000101000000000", -- 513, 512
    513  => "10000000000000000000000000100000001001000000001", -- 514, 513
    514  => "10000000000000000000000000100000001101000000010", -- 515, 514
    515  => "10000000000000000000000000100000010001000000011", -- 516, 515
    516  => "10000000000000000000000000100000010101000000100", -- 517, 516
    517  => "10000000000000000000000000100000011001000000101", -- 518, 517
    518  => "10000000000000000000000000100000011101000000110", -- 519, 518
    519  => "10000000000000000000000000100000100001000000111", -- 520, 519
    520  => "10000000000000000000000000100000100101000001000", -- 521, 520
    521  => "10000000000000000000000000100000101001000001001", -- 522, 521
    522  => "10000000000000000000000000100000101101000001010", -- 523, 522
    523  => "10000000000000000000000000100000110001000001011", -- 524, 523
    524  => "10000000000000000000000000100000110101000001100", -- 525, 524
    525  => "10000000000000000000000000100000111001000001101", -- 526, 525
    526  => "10000000000000000000000000100000111101000001110", -- 527, 526
    527  => "10000000000000000000000000100001000001000001111", -- 528, 527
    528  => "10000000000000000000000000100001000101000010000", -- 529, 528
    529  => "10000000000000000000000000100001001001000010001", -- 530, 529
    530  => "10000000000000000000000000100001001101000010010", -- 531, 530
    531  => "10000000000000000000000000100001010001000010011", -- 532, 531
    532  => "10000000000000000000000000100001010101000010100", -- 533, 532
    533  => "10000000000000000000000000100001011001000010101", -- 534, 533
    534  => "10000000000000000000000000100001011101000010110", -- 535, 534
    535  => "10000000000000000000000000100001100001000010111", -- 536, 535
    536  => "10000000000000000000000000100001100101000011000", -- 537, 536
    537  => "10000000000000000000000000100001101001000011001", -- 538, 537
    538  => "10000000000000000000000000100001101101000011010", -- 539, 538
    539  => "10000000000000000000000000100001110001000011011", -- 540, 539
    540  => "10000000000000000000000000100001110101000011100", -- 541, 540
    541  => "10000000000000000000000000100001111001000011101", -- 542, 541
    542  => "10000000000000000000000000100001111101000011110", -- 543, 542
    543  => "10000000000000000000000000100010000001000011111", -- 544, 543
    544  => "10000000000000000000000000100010000101000100000", -- 545, 544
    545  => "10000000000000000000000000100010001001000100001", -- 546, 545
    546  => "10000000000000000000000000100010001101000100010", -- 547, 546
    547  => "10000000000000000000000000100010010001000100011", -- 548, 547
    548  => "10000000000000000000000000100010010101000100100", -- 549, 548
    549  => "10000000000000000000000000100010011001000100101", -- 550, 549
    550  => "10000000000000000000000000100010011101000100110", -- 551, 550
    551  => "10000000000000000000000000100010100001000100111", -- 552, 551
    552  => "10000000000000000000000000100010100101000101000", -- 553, 552
    553  => "10000000000000000000000000100010101001000101001", -- 554, 553
    554  => "10000000000000000000000000100010101101000101010", -- 555, 554
    555  => "10000000000000000000000000100010110001000101011", -- 556, 555
    556  => "10000000000000000000000000100010110101000101100", -- 557, 556
    557  => "10000000000000000000000000100010111001000101101", -- 558, 557
    558  => "10000000000000000000000000100010111101000101110", -- 559, 558
    559  => "10000000000000000000000000100011000001000101111", -- 560, 559
    560  => "10000000000000000000000000100011000101000110000", -- 561, 560
    561  => "10000000000000000000000000100011001001000110001", -- 562, 561
    562  => "10000000000000000000000000100011001101000110010", -- 563, 562
    563  => "10000000000000000000000000100011010001000110011", -- 564, 563
    564  => "10000000000000000000000000100011010101000110100", -- 565, 564
    565  => "10000000000000000000000000100011011001000110101", -- 566, 565
    566  => "10000000000000000000000000100011011101000110110", -- 567, 566
    567  => "10000000000000000000000000100011100001000110111", -- 568, 567
    568  => "10000000000000000000000000100011100101000111000", -- 569, 568
    569  => "10000000000000000000000000100011101001000111001", -- 570, 569
    570  => "10000000000000000000000000100011101101000111010", -- 571, 570
    571  => "10000000000000000000000000100011110001000111011", -- 572, 571
    572  => "10000000000000000000000000100011110101000111100", -- 573, 572
    573  => "10000000000000000000000000100011111001000111101", -- 574, 573
    574  => "10000000000000000000000000100011111101000111110", -- 575, 574
    575  => "10000000000000000000000000100100000001000111111", -- 576, 575
    576  => "10000000000000000000000000100100000101001000000", -- 577, 576
    577  => "10000000000000000000000000100100001001001000001", -- 578, 577
    578  => "10000000000000000000000000100100001101001000010", -- 579, 578
    579  => "10000000000000000000000000100100010001001000011", -- 580, 579
    580  => "10000000000000000000000000100100010101001000100", -- 581, 580
    581  => "10000000000000000000000000100100011001001000101", -- 582, 581
    582  => "10000000000000000000000000100100011101001000110", -- 583, 582
    583  => "10000000000000000000000000100100100001001000111", -- 584, 583
    584  => "10000000000000000000000000100100100101001001000", -- 585, 584
    585  => "10000000000000000000000000100100101001001001001", -- 586, 585
    586  => "10000000000000000000000000100100101101001001010", -- 587, 586
    587  => "10000000000000000000000000100100110001001001011", -- 588, 587
    588  => "10000000000000000000000000100100110101001001100", -- 589, 588
    589  => "10000000000000000000000000100100111001001001101", -- 590, 589
    590  => "10000000000000000000000000100100111101001001110", -- 591, 590
    591  => "10000000000000000000000000100101000001001001111", -- 592, 591
    592  => "10000000000000000000000000100101000101001010000", -- 593, 592
    593  => "10000000000000000000000000100101001001001010001", -- 594, 593
    594  => "10000000000000000000000000100101001101001010010", -- 595, 594
    595  => "10000000000000000000000000100101010001001010011", -- 596, 595
    596  => "10000000000000000000000000100101010101001010100", -- 597, 596
    597  => "10000000000000000000000000100101011001001010101", -- 598, 597
    598  => "10000000000000000000000000100101011101001010110", -- 599, 598
    599  => "10000000000000000000000000100101100001001010111", -- 600, 599
    600  => "10000000000000000000000000100101100101001011000", -- 601, 600
    601  => "10000000000000000000000000100101101001001011001", -- 602, 601
    602  => "10000000000000000000000000100101101101001011010", -- 603, 602
    603  => "10000000000000000000000000100101110001001011011", -- 604, 603
    604  => "10000000000000000000000000100101110101001011100", -- 605, 604
    605  => "10000000000000000000000000100101111001001011101", -- 606, 605
    606  => "10000000000000000000000000100101111101001011110", -- 607, 606
    607  => "10000000000000000000000000100110000001001011111", -- 608, 607
    608  => "10000000000000000000000000100110000101001100000", -- 609, 608
    609  => "10000000000000000000000000100110001001001100001", -- 610, 609
    610  => "10000000000000000000000000100110001101001100010", -- 611, 610
    611  => "10000000000000000000000000100110010001001100011", -- 612, 611
    612  => "10000000000000000000000000100110010101001100100", -- 613, 612
    613  => "10000000000000000000000000100110011001001100101", -- 614, 613
    614  => "10000000000000000000000000100110011101001100110", -- 615, 614
    615  => "10000000000000000000000000100110100001001100111", -- 616, 615
    616  => "10000000000000000000000000100110100101001101000", -- 617, 616
    617  => "10000000000000000000000000100110101001001101001", -- 618, 617
    618  => "10000000000000000000000000100110101101001101010", -- 619, 618
    619  => "10000000000000000000000000100110110001001101011", -- 620, 619
    620  => "10000000000000000000000000100110110101001101100", -- 621, 620
    621  => "10000000000000000000000000100110111001001101101", -- 622, 621
    622  => "10000000000000000000000000100110111101001101110", -- 623, 622
    623  => "10000000000000000000000000100111000001001101111", -- 624, 623
    624  => "10000000000000000000000000100111000101001110000", -- 625, 624
    625  => "10000000000000000000000000100111001001001110001", -- 626, 625
    626  => "10000000000000000000000000100111001101001110010", -- 627, 626
    627  => "10000000000000000000000000100111010001001110011", -- 628, 627
    628  => "10000000000000000000000000100111010101001110100", -- 629, 628
    629  => "10000000000000000000000000100111011001001110101", -- 630, 629
    630  => "10000000000000000000000000100111011101001110110", -- 631, 630
    631  => "10000000000000000000000000100111100001001110111", -- 632, 631
    632  => "10000000000000000000000000100111100101001111000", -- 633, 632
    633  => "10000000000000000000000000100111101001001111001", -- 634, 633
    634  => "10000000000000000000000000100111101101001111010", -- 635, 634
    635  => "10000000000000000000000000100111110001001111011", -- 636, 635
    636  => "10000000000000000000000000100111110101001111100", -- 637, 636
    637  => "10000000000000000000000000100111111001001111101", -- 638, 637
    638  => "10000000000000000000000000100111111101001111110", -- 639, 638
    639  => "10000000000000000000000000101000000001001111111", -- 640, 639
    640  => "10000000000000000000000000101000000101010000000", -- 641, 640
    641  => "10000000000000000000000000101000001001010000001", -- 642, 641
    642  => "10000000000000000000000000101000001101010000010", -- 643, 642
    643  => "10000000000000000000000000101000010001010000011", -- 644, 643
    644  => "10000000000000000000000000101000010101010000100", -- 645, 644
    645  => "10000000000000000000000000101000011001010000101", -- 646, 645
    646  => "10000000000000000000000000101000011101010000110", -- 647, 646
    647  => "10000000000000000000000000101000100001010000111", -- 648, 647
    648  => "10000000000000000000000000101000100101010001000", -- 649, 648
    649  => "10000000000000000000000000101000101001010001001", -- 650, 649
    650  => "10000000000000000000000000101000101101010001010", -- 651, 650
    651  => "10000000000000000000000000101000110001010001011", -- 652, 651
    652  => "10000000000000000000000000101000110101010001100", -- 653, 652
    653  => "10000000000000000000000000101000111001010001101", -- 654, 653
    654  => "10000000000000000000000000101000111101010001110", -- 655, 654
    655  => "10000000000000000000000000101001000001010001111", -- 656, 655
    656  => "10000000000000000000000000101001000101010010000", -- 657, 656
    657  => "10000000000000000000000000101001001001010010001", -- 658, 657
    658  => "10000000000000000000000000101001001101010010010", -- 659, 658
    659  => "10000000000000000000000000101001010001010010011", -- 660, 659
    660  => "10000000000000000000000000101001010101010010100", -- 661, 660
    661  => "10000000000000000000000000101001011001010010101", -- 662, 661
    662  => "10000000000000000000000000101001011101010010110", -- 663, 662
    663  => "10000000000000000000000000101001100001010010111", -- 664, 663
    664  => "10000000000000000000000000101001100101010011000", -- 665, 664
    665  => "10000000000000000000000000101001101001010011001", -- 666, 665
    666  => "10000000000000000000000000101001101101010011010", -- 667, 666
    667  => "10000000000000000000000000101001110001010011011", -- 668, 667
    668  => "10000000000000000000000000101001110101010011100", -- 669, 668
    669  => "10000000000000000000000000101001111001010011101", -- 670, 669
    670  => "10000000000000000000000000101001111101010011110", -- 671, 670
    671  => "10000000000000000000000000101010000001010011111", -- 672, 671
    672  => "10000000000000000000000000101010000101010100000", -- 673, 672
    673  => "10000000000000000000000000101010001001010100001", -- 674, 673
    674  => "10000000000000000000000000101010001101010100010", -- 675, 674
    675  => "10000000000000000000000000101010010001010100011", -- 676, 675
    676  => "10000000000000000000000000101010010101010100100", -- 677, 676
    677  => "10000000000000000000000000101010011001010100101", -- 678, 677
    678  => "10000000000000000000000000101010011101010100110", -- 679, 678
    679  => "10000000000000000000000000101010100001010100111", -- 680, 679
    680  => "10000000000000000000000000101010100101010101000", -- 681, 680
    681  => "10000000000000000000000000101010101001010101001", -- 682, 681
    682  => "10000000000000000000000000101010101101010101010", -- 683, 682
    683  => "10000000000000000000000000101010110001010101011", -- 684, 683
    684  => "10000000000000000000000000101010110101010101100", -- 685, 684
    685  => "10000000000000000000000000101010111001010101101", -- 686, 685
    686  => "10000000000000000000000000101010111101010101110", -- 687, 686
    687  => "10000000000000000000000000101011000001010101111", -- 688, 687
    688  => "10000000000000000000000000101011000101010110000", -- 689, 688
    689  => "10000000000000000000000000101011001001010110001", -- 690, 689
    690  => "10000000000000000000000000101011001101010110010", -- 691, 690
    691  => "10000000000000000000000000101011010001010110011", -- 692, 691
    692  => "10000000000000000000000000101011010101010110100", -- 693, 692
    693  => "10000000000000000000000000101011011001010110101", -- 694, 693
    694  => "10000000000000000000000000101011011101010110110", -- 695, 694
    695  => "10000000000000000000000000101011100001010110111", -- 696, 695
    696  => "10000000000000000000000000101011100101010111000", -- 697, 696
    697  => "10000000000000000000000000101011101001010111001", -- 698, 697
    698  => "10000000000000000000000000101011101101010111010", -- 699, 698
    699  => "10000000000000000000000000101011110001010111011", -- 700, 699
    700  => "10000000000000000000000000101011110101010111100", -- 701, 700
    701  => "10000000000000000000000000101011111001010111101", -- 702, 701
    702  => "10000000000000000000000000101011111101010111110", -- 703, 702
    703  => "10000000000000000000000000101100000001010111111", -- 704, 703
    704  => "10000000000000000000000000101100000101011000000", -- 705, 704
    705  => "10000000000000000000000000101100001001011000001", -- 706, 705
    706  => "10000000000000000000000000101100001101011000010", -- 707, 706
    707  => "10000000000000000000000000101100010001011000011", -- 708, 707
    708  => "10000000000000000000000000101100010101011000100", -- 709, 708
    709  => "10000000000000000000000000101100011001011000101", -- 710, 709
    710  => "10000000000000000000000000101100011101011000110", -- 711, 710
    711  => "10000000000000000000000000101100100001011000111", -- 712, 711
    712  => "10000000000000000000000000101100100101011001000", -- 713, 712
    713  => "10000000000000000000000000101100101001011001001", -- 714, 713
    714  => "10000000000000000000000000101100101101011001010", -- 715, 714
    715  => "10000000000000000000000000101100110001011001011", -- 716, 715
    716  => "10000000000000000000000000101100110101011001100", -- 717, 716
    717  => "10000000000000000000000000101100111001011001101", -- 718, 717
    718  => "10000000000000000000000000101100111101011001110", -- 719, 718
    719  => "10000000000000000000000000101101000001011001111", -- 720, 719
    720  => "10000000000000000000000000101101000101011010000", -- 721, 720
    721  => "10000000000000000000000000101101001001011010001", -- 722, 721
    722  => "10000000000000000000000000101101001101011010010", -- 723, 722
    723  => "10000000000000000000000000101101010001011010011", -- 724, 723
    724  => "10000000000000000000000000101101010101011010100", -- 725, 724
    725  => "10000000000000000000000000101101011001011010101", -- 726, 725
    726  => "10000000000000000000000000101101011101011010110", -- 727, 726
    727  => "10000000000000000000000000101101100001011010111", -- 728, 727
    728  => "10000000000000000000000000101101100101011011000", -- 729, 728
    729  => "10000000000000000000000000101101101001011011001", -- 730, 729
    730  => "10000000000000000000000000101101101101011011010", -- 731, 730
    731  => "10000000000000000000000000101101110001011011011", -- 732, 731
    732  => "10000000000000000000000000101101110101011011100", -- 733, 732
    733  => "10000000000000000000000000101101111001011011101", -- 734, 733
    734  => "10000000000000000000000000101101111101011011110", -- 735, 734
    735  => "10000000000000000000000000101110000001011011111", -- 736, 735
    736  => "10000000000000000000000000101110000101011100000", -- 737, 736
    737  => "10000000000000000000000000101110001001011100001", -- 738, 737
    738  => "10000000000000000000000000101110001101011100010", -- 739, 738
    739  => "10000000000000000000000000101110010001011100011", -- 740, 739
    740  => "10000000000000000000000000101110010101011100100", -- 741, 740
    741  => "10000000000000000000000000101110011001011100101", -- 742, 741
    742  => "10000000000000000000000000101110011101011100110", -- 743, 742
    743  => "10000000000000000000000000101110100001011100111", -- 744, 743
    744  => "10000000000000000000000000101110100101011101000", -- 745, 744
    745  => "10000000000000000000000000101110101001011101001", -- 746, 745
    746  => "10000000000000000000000000101110101101011101010", -- 747, 746
    747  => "10000000000000000000000000101110110001011101011", -- 748, 747
    748  => "10000000000000000000000000101110110101011101100", -- 749, 748
    749  => "10000000000000000000000000101110111001011101101", -- 750, 749
    750  => "10000000000000000000000000101110111101011101110", -- 751, 750
    751  => "10000000000000000000000000101111000001011101111", -- 752, 751
    752  => "10000000000000000000000000101111000101011110000", -- 753, 752
    753  => "10000000000000000000000000101111001001011110001", -- 754, 753
    754  => "10000000000000000000000000101111001101011110010", -- 755, 754
    755  => "10000000000000000000000000101111010001011110011", -- 756, 755
    756  => "10000000000000000000000000101111010101011110100", -- 757, 756
    757  => "10000000000000000000000000101111011001011110101", -- 758, 757
    758  => "10000000000000000000000000101111011101011110110", -- 759, 758
    759  => "10000000000000000000000000101111100001011110111", -- 760, 759
    760  => "10000000000000000000000000101111100101011111000", -- 761, 760
    761  => "10000000000000000000000000101111101001011111001", -- 762, 761
    762  => "10000000000000000000000000101111101101011111010", -- 763, 762
    763  => "10000000000000000000000000101111110001011111011", -- 764, 763
    764  => "10000000000000000000000000101111110101011111100", -- 765, 764
    765  => "10000000000000000000000000101111111001011111101", -- 766, 765
    766  => "10000000000000000000000000101111111101011111110", -- 767, 766
    767  => "10000000000000000000000000110000000001011111111", -- 768, 767
    768  => "10000000000000000000000000110000000101100000000", -- 769, 768
    769  => "10000000000000000000000000110000001001100000001", -- 770, 769
    770  => "10000000000000000000000000110000001101100000010", -- 771, 770
    771  => "10000000000000000000000000110000010001100000011", -- 772, 771
    772  => "10000000000000000000000000110000010101100000100", -- 773, 772
    773  => "10000000000000000000000000110000011001100000101", -- 774, 773
    774  => "10000000000000000000000000110000011101100000110", -- 775, 774
    775  => "10000000000000000000000000110000100001100000111", -- 776, 775
    776  => "10000000000000000000000000110000100101100001000", -- 777, 776
    777  => "10000000000000000000000000110000101001100001001", -- 778, 777
    778  => "10000000000000000000000000110000101101100001010", -- 779, 778
    779  => "10000000000000000000000000110000110001100001011", -- 780, 779
    780  => "10000000000000000000000000110000110101100001100", -- 781, 780
    781  => "10000000000000000000000000110000111001100001101", -- 782, 781
    782  => "10000000000000000000000000110000111101100001110", -- 783, 782
    783  => "10000000000000000000000000110001000001100001111", -- 784, 783
    784  => "10000000000000000000000000110001000101100010000", -- 785, 784
    785  => "10000000000000000000000000110001001001100010001", -- 786, 785
    786  => "10000000000000000000000000110001001101100010010", -- 787, 786
    787  => "10000000000000000000000000110001010001100010011", -- 788, 787
    788  => "10000000000000000000000000110001010101100010100", -- 789, 788
    789  => "10000000000000000000000000110001011001100010101", -- 790, 789
    790  => "10000000000000000000000000110001011101100010110", -- 791, 790
    791  => "10000000000000000000000000110001100001100010111", -- 792, 791
    792  => "10000000000000000000000000110001100101100011000", -- 793, 792
    793  => "10000000000000000000000000110001101001100011001", -- 794, 793
    794  => "10000000000000000000000000110001101101100011010", -- 795, 794
    795  => "10000000000000000000000000110001110001100011011", -- 796, 795
    796  => "10000000000000000000000000110001110101100011100", -- 797, 796
    797  => "10000000000000000000000000110001111001100011101", -- 798, 797
    798  => "10000000000000000000000000110001111101100011110", -- 799, 798
    799  => "10000000000000000000000000110010000001100011111", -- 800, 799
    800  => "10000000000000000000000000110010000101100100000", -- 801, 800
    801  => "10000000000000000000000000110010001001100100001", -- 802, 801
    802  => "10000000000000000000000000110010001101100100010", -- 803, 802
    803  => "10000000000000000000000000110010010001100100011", -- 804, 803
    804  => "10000000000000000000000000110010010101100100100", -- 805, 804
    805  => "10000000000000000000000000110010011001100100101", -- 806, 805
    806  => "10000000000000000000000000110010011101100100110", -- 807, 806
    807  => "10000000000000000000000000110010100001100100111", -- 808, 807
    808  => "10000000000000000000000000110010100101100101000", -- 809, 808
    809  => "10000000000000000000000000110010101001100101001", -- 810, 809
    810  => "10000000000000000000000000110010101101100101010", -- 811, 810
    811  => "10000000000000000000000000110010110001100101011", -- 812, 811
    812  => "10000000000000000000000000110010110101100101100", -- 813, 812
    813  => "10000000000000000000000000110010111001100101101", -- 814, 813
    814  => "10000000000000000000000000110010111101100101110", -- 815, 814
    815  => "10000000000000000000000000110011000001100101111", -- 816, 815
    816  => "10000000000000000000000000110011000101100110000", -- 817, 816
    817  => "10000000000000000000000000110011001001100110001", -- 818, 817
    818  => "10000000000000000000000000110011001101100110010", -- 819, 818
    819  => "10000000000000000000000000110011010001100110011", -- 820, 819
    820  => "10000000000000000000000000110011010101100110100", -- 821, 820
    821  => "10000000000000000000000000110011011001100110101", -- 822, 821
    822  => "10000000000000000000000000110011011101100110110", -- 823, 822
    823  => "10000000000000000000000000110011100001100110111", -- 824, 823
    824  => "10000000000000000000000000110011100101100111000", -- 825, 824
    825  => "10000000000000000000000000110011101001100111001", -- 826, 825
    826  => "10000000000000000000000000110011101101100111010", -- 827, 826
    827  => "10000000000000000000000000110011110001100111011", -- 828, 827
    828  => "10000000000000000000000000110011110101100111100", -- 829, 828
    829  => "10000000000000000000000000110011111001100111101", -- 830, 829
    830  => "10000000000000000000000000110011111101100111110", -- 831, 830
    831  => "10000000000000000000000000110100000001100111111", -- 832, 831
    832  => "10000000000000000000000000110100000101101000000", -- 833, 832
    833  => "10000000000000000000000000110100001001101000001", -- 834, 833
    834  => "10000000000000000000000000110100001101101000010", -- 835, 834
    835  => "10000000000000000000000000110100010001101000011", -- 836, 835
    836  => "10000000000000000000000000110100010101101000100", -- 837, 836
    837  => "10000000000000000000000000110100011001101000101", -- 838, 837
    838  => "10000000000000000000000000110100011101101000110", -- 839, 838
    839  => "10000000000000000000000000110100100001101000111", -- 840, 839
    840  => "10000000000000000000000000110100100101101001000", -- 841, 840
    841  => "10000000000000000000000000110100101001101001001", -- 842, 841
    842  => "10000000000000000000000000110100101101101001010", -- 843, 842
    843  => "10000000000000000000000000110100110001101001011", -- 844, 843
    844  => "10000000000000000000000000110100110101101001100", -- 845, 844
    845  => "10000000000000000000000000110100111001101001101", -- 846, 845
    846  => "10000000000000000000000000110100111101101001110", -- 847, 846
    847  => "10000000000000000000000000110101000001101001111", -- 848, 847
    848  => "10000000000000000000000000110101000101101010000", -- 849, 848
    849  => "10000000000000000000000000110101001001101010001", -- 850, 849
    850  => "10000000000000000000000000110101001101101010010", -- 851, 850
    851  => "10000000000000000000000000110101010001101010011", -- 852, 851
    852  => "10000000000000000000000000110101010101101010100", -- 853, 852
    853  => "10000000000000000000000000110101011001101010101", -- 854, 853
    854  => "10000000000000000000000000110101011101101010110", -- 855, 854
    855  => "10000000000000000000000000110101100001101010111", -- 856, 855
    856  => "10000000000000000000000000110101100101101011000", -- 857, 856
    857  => "10000000000000000000000000110101101001101011001", -- 858, 857
    858  => "10000000000000000000000000110101101101101011010", -- 859, 858
    859  => "10000000000000000000000000110101110001101011011", -- 860, 859
    860  => "10000000000000000000000000110101110101101011100", -- 861, 860
    861  => "10000000000000000000000000110101111001101011101", -- 862, 861
    862  => "10000000000000000000000000110101111101101011110", -- 863, 862
    863  => "10000000000000000000000000110110000001101011111", -- 864, 863
    864  => "10000000000000000000000000110110000101101100000", -- 865, 864
    865  => "10000000000000000000000000110110001001101100001", -- 866, 865
    866  => "10000000000000000000000000110110001101101100010", -- 867, 866
    867  => "10000000000000000000000000110110010001101100011", -- 868, 867
    868  => "10000000000000000000000000110110010101101100100", -- 869, 868
    869  => "10000000000000000000000000110110011001101100101", -- 870, 869
    870  => "10000000000000000000000000110110011101101100110", -- 871, 870
    871  => "10000000000000000000000000110110100001101100111", -- 872, 871
    872  => "10000000000000000000000000110110100101101101000", -- 873, 872
    873  => "10000000000000000000000000110110101001101101001", -- 874, 873
    874  => "10000000000000000000000000110110101101101101010", -- 875, 874
    875  => "10000000000000000000000000110110110001101101011", -- 876, 875
    876  => "10000000000000000000000000110110110101101101100", -- 877, 876
    877  => "10000000000000000000000000110110111001101101101", -- 878, 877
    878  => "10000000000000000000000000110110111101101101110", -- 879, 878
    879  => "10000000000000000000000000110111000001101101111", -- 880, 879
    880  => "10000000000000000000000000110111000101101110000", -- 881, 880
    881  => "10000000000000000000000000110111001001101110001", -- 882, 881
    882  => "10000000000000000000000000110111001101101110010", -- 883, 882
    883  => "10000000000000000000000000110111010001101110011", -- 884, 883
    884  => "10000000000000000000000000110111010101101110100", -- 885, 884
    885  => "10000000000000000000000000110111011001101110101", -- 886, 885
    886  => "10000000000000000000000000110111011101101110110", -- 887, 886
    887  => "10000000000000000000000000110111100001101110111", -- 888, 887
    888  => "10000000000000000000000000110111100101101111000", -- 889, 888
    889  => "10000000000000000000000000110111101001101111001", -- 890, 889
    890  => "10000000000000000000000000110111101101101111010", -- 891, 890
    891  => "10000000000000000000000000110111110001101111011", -- 892, 891
    892  => "10000000000000000000000000110111110101101111100", -- 893, 892
    893  => "10000000000000000000000000110111111001101111101", -- 894, 893
    894  => "10000000000000000000000000110111111101101111110", -- 895, 894
    895  => "10000000000000000000000000111000000001101111111", -- 896, 895
    896  => "10000000000000000000000000111000000101110000000", -- 897, 896
    897  => "10000000000000000000000000111000001001110000001", -- 898, 897
    898  => "10000000000000000000000000111000001101110000010", -- 899, 898
    899  => "10000000000000000000000000111000010001110000011", -- 900, 899
    900  => "10000000000000000000000000111000010101110000100", -- 901, 900
    901  => "10000000000000000000000000111000011001110000101", -- 902, 901
    902  => "10000000000000000000000000111000011101110000110", -- 903, 902
    903  => "10000000000000000000000000111000100001110000111", -- 904, 903
    904  => "10000000000000000000000000111000100101110001000", -- 905, 904
    905  => "10000000000000000000000000111000101001110001001", -- 906, 905
    906  => "10000000000000000000000000111000101101110001010", -- 907, 906
    907  => "10000000000000000000000000111000110001110001011", -- 908, 907
    908  => "10000000000000000000000000111000110101110001100", -- 909, 908
    909  => "10000000000000000000000000111000111001110001101", -- 910, 909
    910  => "10000000000000000000000000111000111101110001110", -- 911, 910
    911  => "10000000000000000000000000111001000001110001111", -- 912, 911
    912  => "10000000000000000000000000111001000101110010000", -- 913, 912
    913  => "10000000000000000000000000111001001001110010001", -- 914, 913
    914  => "10000000000000000000000000111001001101110010010", -- 915, 914
    915  => "10000000000000000000000000111001010001110010011", -- 916, 915
    916  => "10000000000000000000000000111001010101110010100", -- 917, 916
    917  => "10000000000000000000000000111001011001110010101", -- 918, 917
    918  => "10000000000000000000000000111001011101110010110", -- 919, 918
    919  => "10000000000000000000000000111001100001110010111", -- 920, 919
    920  => "10000000000000000000000000111001100101110011000", -- 921, 920
    921  => "10000000000000000000000000111001101001110011001", -- 922, 921
    922  => "10000000000000000000000000111001101101110011010", -- 923, 922
    923  => "10000000000000000000000000111001110001110011011", -- 924, 923
    924  => "10000000000000000000000000111001110101110011100", -- 925, 924
    925  => "10000000000000000000000000111001111001110011101", -- 926, 925
    926  => "10000000000000000000000000111001111101110011110", -- 927, 926
    927  => "10000000000000000000000000111010000001110011111", -- 928, 927
    928  => "10000000000000000000000000111010000101110100000", -- 929, 928
    929  => "10000000000000000000000000111010001001110100001", -- 930, 929
    930  => "10000000000000000000000000111010001101110100010", -- 931, 930
    931  => "10000000000000000000000000111010010001110100011", -- 932, 931
    932  => "10000000000000000000000000111010010101110100100", -- 933, 932
    933  => "10000000000000000000000000111010011001110100101", -- 934, 933
    934  => "10000000000000000000000000111010011101110100110", -- 935, 934
    935  => "10000000000000000000000000111010100001110100111", -- 936, 935
    936  => "10000000000000000000000000111010100101110101000", -- 937, 936
    937  => "10000000000000000000000000111010101001110101001", -- 938, 937
    938  => "10000000000000000000000000111010101101110101010", -- 939, 938
    939  => "10000000000000000000000000111010110001110101011", -- 940, 939
    940  => "10000000000000000000000000111010110101110101100", -- 941, 940
    941  => "10000000000000000000000000111010111001110101101", -- 942, 941
    942  => "10000000000000000000000000111010111101110101110", -- 943, 942
    943  => "10000000000000000000000000111011000001110101111", -- 944, 943
    944  => "10000000000000000000000000111011000101110110000", -- 945, 944
    945  => "10000000000000000000000000111011001001110110001", -- 946, 945
    946  => "10000000000000000000000000111011001101110110010", -- 947, 946
    947  => "10000000000000000000000000111011010001110110011", -- 948, 947
    948  => "10000000000000000000000000111011010101110110100", -- 949, 948
    949  => "10000000000000000000000000111011011001110110101", -- 950, 949
    950  => "10000000000000000000000000111011011101110110110", -- 951, 950
    951  => "10000000000000000000000000111011100001110110111", -- 952, 951
    952  => "10000000000000000000000000111011100101110111000", -- 953, 952
    953  => "10000000000000000000000000111011101001110111001", -- 954, 953
    954  => "10000000000000000000000000111011101101110111010", -- 955, 954
    955  => "10000000000000000000000000111011110001110111011", -- 956, 955
    956  => "10000000000000000000000000111011110101110111100", -- 957, 956
    957  => "10000000000000000000000000111011111001110111101", -- 958, 957
    958  => "10000000000000000000000000111011111101110111110", -- 959, 958
    959  => "10000000000000000000000000111100000001110111111", -- 960, 959
    960  => "10000000000000000000000000111100000101111000000", -- 961, 960
    961  => "10000000000000000000000000111100001001111000001", -- 962, 961
    962  => "10000000000000000000000000111100001101111000010", -- 963, 962
    963  => "10000000000000000000000000111100010001111000011", -- 964, 963
    964  => "10000000000000000000000000111100010101111000100", -- 965, 964
    965  => "10000000000000000000000000111100011001111000101", -- 966, 965
    966  => "10000000000000000000000000111100011101111000110", -- 967, 966
    967  => "10000000000000000000000000111100100001111000111", -- 968, 967
    968  => "10000000000000000000000000111100100101111001000", -- 969, 968
    969  => "10000000000000000000000000111100101001111001001", -- 970, 969
    970  => "10000000000000000000000000111100101101111001010", -- 971, 970
    971  => "10000000000000000000000000111100110001111001011", -- 972, 971
    972  => "10000000000000000000000000111100110101111001100", -- 973, 972
    973  => "10000000000000000000000000111100111001111001101", -- 974, 973
    974  => "10000000000000000000000000111100111101111001110", -- 975, 974
    975  => "10000000000000000000000000111101000001111001111", -- 976, 975
    976  => "10000000000000000000000000111101000101111010000", -- 977, 976
    977  => "10000000000000000000000000111101001001111010001", -- 978, 977
    978  => "10000000000000000000000000111101001101111010010", -- 979, 978
    979  => "10000000000000000000000000111101010001111010011", -- 980, 979
    980  => "10000000000000000000000000111101010101111010100", -- 981, 980
    981  => "10000000000000000000000000111101011001111010101", -- 982, 981
    982  => "10000000000000000000000000111101011101111010110", -- 983, 982
    983  => "10000000000000000000000000111101100001111010111", -- 984, 983
    984  => "10000000000000000000000000111101100101111011000", -- 985, 984
    985  => "10000000000000000000000000111101101001111011001", -- 986, 985
    986  => "10000000000000000000000000111101101101111011010", -- 987, 986
    987  => "10000000000000000000000000111101110001111011011", -- 988, 987
    988  => "10000000000000000000000000111101110101111011100", -- 989, 988
    989  => "10000000000000000000000000111101111001111011101", -- 990, 989
    990  => "10000000000000000000000000111101111101111011110", -- 991, 990
    991  => "10000000000000000000000000111110000001111011111", -- 992, 991
    992  => "10000000000000000000000000111110000101111100000", -- 993, 992
    993  => "10000000000000000000000000111110001001111100001", -- 994, 993
    994  => "10000000000000000000000000111110001101111100010", -- 995, 994
    995  => "10000000000000000000000000111110010001111100011", -- 996, 995
    996  => "10000000000000000000000000111110010101111100100", -- 997, 996
    997  => "10000000000000000000000000111110011001111100101", -- 998, 997
    998  => "10000000000000000000000000111110011101111100110", -- 999, 998
    999  => "10000000000000000000000000111110100001111100111", -- 1000, 999
    1000 => "10000000000000000000000000111110100101111101000", -- 1001, 1000
    1001 => "10000000000000000000000000111110101001111101001", -- 1002, 1001
    1002 => "10000000000000000000000000111110101101111101010", -- 1003, 1002
    1003 => "10000000000000000000000000111110110001111101011", -- 1004, 1003
    1004 => "10000000000000000000000000111110110101111101100", -- 1005, 1004
    1005 => "10000000000000000000000000111110111001111101101", -- 1006, 1005
    1006 => "10000000000000000000000000111110111101111101110", -- 1007, 1006
    1007 => "10000000000000000000000000111111000001111101111", -- 1008, 1007
    1008 => "10000000000000000000000000111111000101111110000", -- 1009, 1008
    1009 => "10000000000000000000000000111111001001111110001", -- 1010, 1009
    1010 => "10000000000000000000000000111111001101111110010", -- 1011, 1010
    1011 => "10000000000000000000000000111111010001111110011", -- 1012, 1011
    1012 => "10000000000000000000000000111111010101111110100", -- 1013, 1012
    1013 => "10000000000000000000000000111111011001111110101", -- 1014, 1013
    1014 => "10000000000000000000000000111111011101111110110", -- 1015, 1014
    1015 => "10000000000000000000000000111111100001111110111", -- 1016, 1015
    1016 => "10000000000000000000000000111111100101111111000", -- 1017, 1016
    1017 => "10000000000000000000000000111111101001111111001", -- 1018, 1017
    1018 => "10000000000000000000000000111111101101111111010", -- 1019, 1018
    1019 => "10000000000000000000000000111111110001111111011", -- 1020, 1019
    1020 => "10000000000000000000000000111111110101111111100", -- 1021, 1020
    1021 => "10000000000000000000000000111111111001111111101", -- 1022, 1021
    1022 => "10000000000000000000000000111111111101111111110", -- 1023, 1022
    1023 => "10000000000000000000000001111111111101111111111" -- null, 1023
  );

  constant init_rate_mem_1024 : rate_mem_type := (
    0    => "001101001",
    1    => "110110000",
    2    => "100000001",
    3    => "110000111",
    4    => "001111010",
    5    => "010001111",
    6    => "101010001",
    7    => "001001001",
    8    => "110111010",
    9    => "000101011",
    10   => "011010110",
    11   => "111000000",
    12   => "101011010",
    13   => "010001000",
    14   => "101101101",
    15   => "100101111",
    16   => "000010001",
    17   => "100001010",
    18   => "110110010",
    19   => "111011010",
    20   => "111011100",
    21   => "011110001",
    22   => "010110100",
    23   => "101101101",
    24   => "010000100",
    25   => "001010100",
    26   => "000010101",
    27   => "100000111",
    28   => "111001100",
    29   => "110111000",
    30   => "010101111",
    31   => "011010000",
    32   => "011110110",
    33   => "010100000",
    34   => "010011101",
    35   => "000111001",
    36   => "011011111",
    37   => "000010010",
    38   => "001001011",
    39   => "011000101",
    40   => "001000000",
    41   => "110110000",
    42   => "001100010",
    43   => "000111111",
    44   => "110001010",
    45   => "110111110",
    46   => "110011011",
    47   => "001100110",
    48   => "100111101",
    49   => "001010011",
    50   => "001101010",
    51   => "010011101",
    52   => "111010111",
    53   => "011001000",
    54   => "011000110",
    55   => "100010100",
    56   => "111001100",
    57   => "001100110",
    58   => "000100011",
    59   => "011111110",
    60   => "011111000",
    61   => "010010000",
    62   => "111000101",
    63   => "110101100",
    64   => "101110001",
    65   => "010110100",
    66   => "111101110",
    67   => "010010101",
    68   => "010101111",
    69   => "101011011",
    70   => "001110111",
    71   => "100000011",
    72   => "100010000",
    73   => "111101100",
    74   => "001111011",
    75   => "110111100",
    76   => "001010101",
    77   => "011100100",
    78   => "011000011",
    79   => "011110001",
    80   => "000010000",
    81   => "110011001",
    82   => "111011011",
    83   => "001100011",
    84   => "100101110",
    85   => "111111001",
    86   => "101100111",
    87   => "011011110",
    88   => "111010111",
    89   => "010111100",
    90   => "010010000",
    91   => "010100010",
    92   => "011000010",
    93   => "100110010",
    94   => "100000010",
    95   => "000101101",
    96   => "010100010",
    97   => "111111010",
    98   => "000010011",
    99   => "011011011",
    100  => "111100100",
    101  => "100110000",
    102  => "101000010",
    103  => "001001001",
    104  => "110101110",
    105  => "010001100",
    106  => "101011100",
    107  => "100110111",
    108  => "101100001",
    109  => "011000111",
    110  => "011011111",
    111  => "110111011",
    112  => "101010111",
    113  => "110001011",
    114  => "001001011",
    115  => "110111011",
    116  => "110000100",
    117  => "011000000",
    118  => "001011100",
    119  => "010100110",
    120  => "111101110",
    121  => "000011100",
    122  => "100011110",
    123  => "110111111",
    124  => "001000101",
    125  => "110000010",
    126  => "111111110",
    127  => "110101110",
    128  => "010100001",
    129  => "001000100",
    130  => "100110000",
    131  => "001001101",
    132  => "111010110",
    133  => "000110101",
    134  => "110001001",
    135  => "101000000",
    136  => "011111111",
    137  => "011110100",
    138  => "100010011",
    139  => "101100000",
    140  => "010100101",
    141  => "010011100",
    142  => "010011011",
    143  => "110111000",
    144  => "111100111",
    145  => "001110111",
    146  => "110011100",
    147  => "000001100",
    148  => "001110110",
    149  => "010101011",
    150  => "100011101",
    151  => "001110011",
    152  => "101110011",
    153  => "011001001",
    154  => "110001101",
    155  => "010001000",
    156  => "111100110",
    157  => "100110101",
    158  => "010000000",
    159  => "001001100",
    160  => "100011110",
    161  => "101100000",
    162  => "001010011",
    163  => "101100101",
    164  => "011011001",
    165  => "100011111",
    166  => "110001101",
    167  => "011101101",
    168  => "110001011",
    169  => "001000010",
    170  => "101011110",
    171  => "010100000",
    172  => "010001101",
    173  => "110010011",
    174  => "111001011",
    175  => "000010111",
    176  => "110010000",
    177  => "100010111",
    178  => "111111111",
    179  => "101111111",
    180  => "001001011",
    181  => "010100010",
    182  => "101111101",
    183  => "110011001",
    184  => "000110001",
    185  => "001000100",
    186  => "101000000",
    187  => "110101100",
    188  => "001110101",
    189  => "101101001",
    190  => "100010111",
    191  => "001101100",
    192  => "100101101",
    193  => "010010011",
    194  => "101101100",
    195  => "001000111",
    196  => "011001111",
    197  => "101111000",
    198  => "101110100",
    199  => "010101011",
    200  => "011110110",
    201  => "111010101",
    202  => "111001111",
    203  => "001100110",
    204  => "001111101",
    205  => "101110101",
    206  => "100101101",
    207  => "010111100",
    208  => "111100001",
    209  => "010010111",
    210  => "000010101",
    211  => "101110001",
    212  => "110110011",
    213  => "100000001",
    214  => "110101101",
    215  => "100111111",
    216  => "010111111",
    217  => "001101010",
    218  => "000011110",
    219  => "010000111",
    220  => "100100111",
    221  => "101000110",
    222  => "101010010",
    223  => "000001101",
    224  => "010100101",
    225  => "011001010",
    226  => "000001110",
    227  => "111110111",
    228  => "000010110",
    229  => "011101010",
    230  => "111000100",
    231  => "100010001",
    232  => "010011001",
    233  => "001100100",
    234  => "001111011",
    235  => "101011101",
    236  => "001000110",
    237  => "110111101",
    238  => "101001011",
    239  => "101110100",
    240  => "100101111",
    241  => "110111110",
    242  => "010101001",
    243  => "000011100",
    244  => "101111110",
    245  => "010101011",
    246  => "000010100",
    247  => "101010111",
    248  => "110001000",
    249  => "000111011",
    250  => "000100000",
    251  => "100001010",
    252  => "010011011",
    253  => "001000000",
    254  => "011011010",
    255  => "111110001",
    256  => "011011001",
    257  => "100000111",
    258  => "100100101",
    259  => "111010111",
    260  => "001001010",
    261  => "100001101",
    262  => "000111100",
    263  => "110010011",
    264  => "011101000",
    265  => "001000100",
    266  => "000101110",
    267  => "110011000",
    268  => "001111111",
    269  => "011010110",
    270  => "001100010",
    271  => "110110101",
    272  => "111000101",
    273  => "001011111",
    274  => "111110100",
    275  => "000010001",
    276  => "100001011",
    277  => "011100000",
    278  => "000100101",
    279  => "011111010",
    280  => "001110001",
    281  => "011000010",
    282  => "110111111",
    283  => "010111110",
    284  => "011101100",
    285  => "111010100",
    286  => "001000100",
    287  => "111110100",
    288  => "011100100",
    289  => "110001111",
    290  => "100011010",
    291  => "110100111",
    292  => "100100110",
    293  => "011101110",
    294  => "101100000",
    295  => "111110001",
    296  => "011100111",
    297  => "001001110",
    298  => "001000011",
    299  => "111001000",
    300  => "101011100",
    301  => "011111110",
    302  => "111101110",
    303  => "100000001",
    304  => "010101011",
    305  => "010100111",
    306  => "110000011",
    307  => "111011110",
    308  => "000001100",
    309  => "110011010",
    310  => "111100101",
    311  => "111110000",
    312  => "110110100",
    313  => "110101111",
    314  => "110000010",
    315  => "001111100",
    316  => "110001101",
    317  => "001011010",
    318  => "110101010",
    319  => "001000100",
    320  => "100000110",
    321  => "011011110",
    322  => "100110100",
    323  => "100010000",
    324  => "100101101",
    325  => "000011100",
    326  => "011110110",
    327  => "100101010",
    328  => "010111011",
    329  => "000111101",
    330  => "010001111",
    331  => "011010110",
    332  => "101110100",
    333  => "100000000",
    334  => "001011000",
    335  => "110011001",
    336  => "110010101",
    337  => "011101001",
    338  => "001100000",
    339  => "111101101",
    340  => "011101000",
    341  => "001110100",
    342  => "011111000",
    343  => "000011110",
    344  => "001100010",
    345  => "100010001",
    346  => "111000010",
    347  => "110011000",
    348  => "011110001",
    349  => "110000101",
    350  => "110111111",
    351  => "001010100",
    352  => "010111111",
    353  => "011111011",
    354  => "111101001",
    355  => "101101101",
    356  => "111010010",
    357  => "100101111",
    358  => "110100010",
    359  => "100101001",
    360  => "101101100",
    361  => "110000111",
    362  => "001110000",
    363  => "101011110",
    364  => "111000010",
    365  => "110001111",
    366  => "101101010",
    367  => "001000100",
    368  => "011010010",
    369  => "011011010",
    370  => "111110110",
    371  => "000110010",
    372  => "011011000",
    373  => "110100110",
    374  => "000111111",
    375  => "100011000",
    376  => "011101011",
    377  => "110111110",
    378  => "010001001",
    379  => "001101111",
    380  => "010110001",
    381  => "100100101",
    382  => "110111101",
    383  => "111010000",
    384  => "110100101",
    385  => "000111100",
    386  => "001011011",
    387  => "010000111",
    388  => "001010110",
    389  => "001101110",
    390  => "110100000",
    391  => "100010111",
    392  => "100101101",
    393  => "101000100",
    394  => "101010010",
    395  => "111111100",
    396  => "010111101",
    397  => "101111110",
    398  => "100110010",
    399  => "011010010",
    400  => "010001001",
    401  => "011000111",
    402  => "000111010",
    403  => "101011101",
    404  => "100100011",
    405  => "011011111",
    406  => "010010001",
    407  => "100000000",
    408  => "000101010",
    409  => "110110000",
    410  => "101010110",
    411  => "111011011",
    412  => "101101001",
    413  => "110011000",
    414  => "010010100",
    415  => "111100011",
    416  => "100110110",
    417  => "000001111",
    418  => "101001001",
    419  => "000101010",
    420  => "101000001",
    421  => "001000100",
    422  => "111111001",
    423  => "111111110",
    424  => "111110001",
    425  => "100011101",
    426  => "011111110",
    427  => "001100100",
    428  => "110010001",
    429  => "001000110",
    430  => "111110100",
    431  => "000111000",
    432  => "010100100",
    433  => "010100101",
    434  => "101101101",
    435  => "111001011",
    436  => "101111001",
    437  => "001000110",
    438  => "001000101",
    439  => "011110110",
    440  => "011011110",
    441  => "101101010",
    442  => "111010010",
    443  => "000101001",
    444  => "100011000",
    445  => "001100001",
    446  => "111001010",
    447  => "110100011",
    448  => "010011111",
    449  => "011011100",
    450  => "001100101",
    451  => "100011001",
    452  => "010101011",
    453  => "001011011",
    454  => "000111100",
    455  => "011011110",
    456  => "000100011",
    457  => "100111010",
    458  => "011000100",
    459  => "011011011",
    460  => "100010100",
    461  => "011001100",
    462  => "000111000",
    463  => "010000111",
    464  => "100000101",
    465  => "110100101",
    466  => "110101011",
    467  => "111110011",
    468  => "001000011",
    469  => "011011110",
    470  => "010001101",
    471  => "000110000",
    472  => "011010101",
    473  => "111001010",
    474  => "101010000",
    475  => "001001001",
    476  => "000010000",
    477  => "011001100",
    478  => "000001101",
    479  => "000001110",
    480  => "111111100",
    481  => "111101000",
    482  => "001010001",
    483  => "101001110",
    484  => "100001011",
    485  => "111000011",
    486  => "111101111",
    487  => "000101101",
    488  => "011001001",
    489  => "001000000",
    490  => "001011001",
    491  => "011001011",
    492  => "101000111",
    493  => "100110000",
    494  => "001110111",
    495  => "111010110",
    496  => "011011001",
    497  => "000111000",
    498  => "101111100",
    499  => "110001111",
    500  => "011111000",
    501  => "100100100",
    502  => "101110101",
    503  => "101111100",
    504  => "101101001",
    505  => "111000000",
    506  => "010111111",
    507  => "100011100",
    508  => "101001101",
    509  => "000011110",
    510  => "000101101",
    511  => "111010101",
    512  => "100101100",
    513  => "010010011",
    514  => "000011110",
    515  => "011000011",
    516  => "101100010",
    517  => "011011101",
    518  => "010100010",
    519  => "010111010",
    520  => "010111101",
    521  => "111011100",
    522  => "111100101",
    523  => "001101100",
    524  => "101100001",
    525  => "100111000",
    526  => "110101111",
    527  => "000110111",
    528  => "101111100",
    529  => "101011010",
    530  => "100101110",
    531  => "100001010",
    532  => "111101111",
    533  => "000001101",
    534  => "001000111",
    535  => "111101101",
    536  => "011000011",
    537  => "000001101",
    538  => "111001010",
    539  => "110100100",
    540  => "110101000",
    541  => "010101010",
    542  => "000100110",
    543  => "101111110",
    544  => "110000100",
    545  => "101110010",
    546  => "010110100",
    547  => "110000111",
    548  => "101111111",
    549  => "010100010",
    550  => "110001111",
    551  => "101101001",
    552  => "011010000",
    553  => "111100010",
    554  => "000011010",
    555  => "011110000",
    556  => "100111101",
    557  => "001011001",
    558  => "101111001",
    559  => "001101111",
    560  => "110100111",
    561  => "111110111",
    562  => "000110011",
    563  => "110110011",
    564  => "010011101",
    565  => "110000101",
    566  => "101111010",
    567  => "001100010",
    568  => "110110010",
    569  => "101110011",
    570  => "100101011",
    571  => "100000001",
    572  => "010111011",
    573  => "111111101",
    574  => "111010001",
    575  => "110111100",
    576  => "000111010",
    577  => "011110111",
    578  => "010010111",
    579  => "011001010",
    580  => "101011010",
    581  => "111001100",
    582  => "010001011",
    583  => "011100011",
    584  => "110000000",
    585  => "010111110",
    586  => "011110010",
    587  => "101100101",
    588  => "001010101",
    589  => "110110101",
    590  => "011000100",
    591  => "110001011",
    592  => "010111000",
    593  => "101000000",
    594  => "100111011",
    595  => "011110011",
    596  => "010101111",
    597  => "001100101",
    598  => "010000110",
    599  => "101000101",
    600  => "110100100",
    601  => "110101101",
    602  => "011000010",
    603  => "111001111",
    604  => "100110100",
    605  => "011011011",
    606  => "010111100",
    607  => "000011010",
    608  => "010101010",
    609  => "111110011",
    610  => "001110000",
    611  => "010001100",
    612  => "010111111",
    613  => "001100101",
    614  => "010100101",
    615  => "111000011",
    616  => "100000100",
    617  => "001101000",
    618  => "001001000",
    619  => "001001100",
    620  => "011010000",
    621  => "010001111",
    622  => "000100000",
    623  => "010001010",
    624  => "000011001",
    625  => "111101011",
    626  => "111100100",
    627  => "010100000",
    628  => "110011010",
    629  => "010110101",
    630  => "001100100",
    631  => "111000011",
    632  => "111001110",
    633  => "110111000",
    634  => "101101100",
    635  => "000100101",
    636  => "110100000",
    637  => "111000101",
    638  => "110111100",
    639  => "101100110",
    640  => "010110111",
    641  => "110100000",
    642  => "110010100",
    643  => "111101100",
    644  => "100111101",
    645  => "111111011",
    646  => "011001100",
    647  => "100000000",
    648  => "110010110",
    649  => "001000000",
    650  => "000011101",
    651  => "011000000",
    652  => "110111011",
    653  => "000011000",
    654  => "000111011",
    655  => "010001010",
    656  => "111110001",
    657  => "011100011",
    658  => "110001001",
    659  => "110010110",
    660  => "100100001",
    661  => "011001100",
    662  => "001011110",
    663  => "000110111",
    664  => "101111011",
    665  => "100010000",
    666  => "111100011",
    667  => "001001111",
    668  => "001001010",
    669  => "011011101",
    670  => "110100000",
    671  => "010101001",
    672  => "010110010",
    673  => "010001101",
    674  => "111100000",
    675  => "101111000",
    676  => "011110111",
    677  => "100100011",
    678  => "100101000",
    679  => "111110100",
    680  => "001101000",
    681  => "010100111",
    682  => "001001010",
    683  => "000111110",
    684  => "111100011",
    685  => "000100111",
    686  => "110101110",
    687  => "101111110",
    688  => "001010011",
    689  => "101011001",
    690  => "110000011",
    691  => "010001001",
    692  => "110001111",
    693  => "011101010",
    694  => "001100110",
    695  => "110010110",
    696  => "001101110",
    697  => "110010001",
    698  => "010110001",
    699  => "001111011",
    700  => "000001011",
    701  => "011111110",
    702  => "111011111",
    703  => "101001101",
    704  => "100000000",
    705  => "110101001",
    706  => "100010000",
    707  => "101010100",
    708  => "001000100",
    709  => "110001010",
    710  => "010111011",
    711  => "001100100",
    712  => "110100110",
    713  => "011101111",
    714  => "111110101",
    715  => "111110100",
    716  => "010000001",
    717  => "101000001",
    718  => "100101011",
    719  => "100111101",
    720  => "000010010",
    721  => "101011101",
    722  => "001000011",
    723  => "100111110",
    724  => "011010101",
    725  => "011101101",
    726  => "011000111",
    727  => "001010111",
    728  => "110001010",
    729  => "110000100",
    730  => "001111100",
    731  => "010010100",
    732  => "100110110",
    733  => "010110111",
    734  => "101100101",
    735  => "010000110",
    736  => "111110000",
    737  => "001101110",
    738  => "011100101",
    739  => "000111010",
    740  => "101110011",
    741  => "111011010",
    742  => "010100000",
    743  => "011011000",
    744  => "001111111",
    745  => "010110000",
    746  => "011111101",
    747  => "010111101",
    748  => "011100100",
    749  => "101111111",
    750  => "001111100",
    751  => "101100101",
    752  => "110111001",
    753  => "101110111",
    754  => "100000111",
    755  => "110100000",
    756  => "101100011",
    757  => "101100011",
    758  => "001101101",
    759  => "111000111",
    760  => "001001110",
    761  => "111010111",
    762  => "001111001",
    763  => "010011001",
    764  => "011011011",
    765  => "010111111",
    766  => "001101010",
    767  => "111010101",
    768  => "100000000",
    769  => "010110001",
    770  => "000010100",
    771  => "001001010",
    772  => "111111000",
    773  => "100001101",
    774  => "011010100",
    775  => "100101001",
    776  => "101100111",
    777  => "011111101",
    778  => "101111110",
    779  => "111100010",
    780  => "100000110",
    781  => "111011110",
    782  => "010011010",
    783  => "111101000",
    784  => "111000110",
    785  => "110101100",
    786  => "110001111",
    787  => "011000111",
    788  => "100101001",
    789  => "000101100",
    790  => "101000000",
    791  => "100101110",
    792  => "001110101",
    793  => "000010001",
    794  => "101010100",
    795  => "111000000",
    796  => "010100000",
    797  => "100111000",
    798  => "001111101",
    799  => "011011010",
    800  => "110001110",
    801  => "100000000",
    802  => "000001110",
    803  => "100111011",
    804  => "111110010",
    805  => "110010011",
    806  => "110001100",
    807  => "001010010",
    808  => "110100110",
    809  => "100001000",
    810  => "001010101",
    811  => "011011100",
    812  => "001000100",
    813  => "111111000",
    814  => "011001110",
    815  => "001011001",
    816  => "101011110",
    817  => "111010111",
    818  => "111111111",
    819  => "111110101",
    820  => "001110111",
    821  => "110110001",
    822  => "000010011",
    823  => "111111111",
    824  => "001101111",
    825  => "111101011",
    826  => "011110011",
    827  => "101010101",
    828  => "011100111",
    829  => "011011101",
    830  => "001010110",
    831  => "111001110",
    832  => "100110100",
    833  => "110001011",
    834  => "101010111",
    835  => "111011101",
    836  => "111001010",
    837  => "110100100",
    838  => "101110111",
    839  => "110010110",
    840  => "011101101",
    841  => "101010010",
    842  => "000101111",
    843  => "010000010",
    844  => "110010001",
    845  => "011000011",
    846  => "011011100",
    847  => "010010111",
    848  => "001010100",
    849  => "101100101",
    850  => "101101111",
    851  => "000101011",
    852  => "000101110",
    853  => "001010011",
    854  => "111100101",
    855  => "110110011",
    856  => "011101110",
    857  => "000101111",
    858  => "100000111",
    859  => "000101110",
    860  => "110101011",
    861  => "001000111",
    862  => "100110010",
    863  => "111111101",
    864  => "010110001",
    865  => "100011010",
    866  => "011010101",
    867  => "100010101",
    868  => "001111000",
    869  => "010110101",
    870  => "000011111",
    871  => "101011111",
    872  => "111001101",
    873  => "110001011",
    874  => "011010101",
    875  => "110111100",
    876  => "110101100",
    877  => "111110010",
    878  => "001010100",
    879  => "110100110",
    880  => "010100111",
    881  => "101110001",
    882  => "011010110",
    883  => "101111111",
    884  => "001101010",
    885  => "010011110",
    886  => "111010011",
    887  => "101101010",
    888  => "000110110",
    889  => "011111011",
    890  => "111110000",
    891  => "111111101",
    892  => "001110001",
    893  => "111111101",
    894  => "000011000",
    895  => "010100111",
    896  => "101001010",
    897  => "100001000",
    898  => "011101111",
    899  => "000100001",
    900  => "011000110",
    901  => "100100101",
    902  => "100110011",
    903  => "010001010",
    904  => "100100111",
    905  => "001111011",
    906  => "100100101",
    907  => "110010000",
    908  => "110100011",
    909  => "000110110",
    910  => "110110101",
    911  => "100100010",
    912  => "101101111",
    913  => "001001011",
    914  => "000101111",
    915  => "101110100",
    916  => "101001100",
    917  => "011000111",
    918  => "011111100",
    919  => "001011110",
    920  => "001111010",
    921  => "101011100",
    922  => "010010110",
    923  => "011101011",
    924  => "001111011",
    925  => "001110100",
    926  => "010001011",
    927  => "010111101",
    928  => "001001101",
    929  => "010010100",
    930  => "010110010",
    931  => "101110000",
    932  => "100111101",
    933  => "001111101",
    934  => "011101010",
    935  => "101001001",
    936  => "110001011",
    937  => "010010110",
    938  => "100001101",
    939  => "100101000",
    940  => "100001011",
    941  => "010000100",
    942  => "011001010",
    943  => "111111001",
    944  => "101111010",
    945  => "100100100",
    946  => "111101101",
    947  => "011011101",
    948  => "010011001",
    949  => "111111111",
    950  => "111110111",
    951  => "011111111",
    952  => "011011101",
    953  => "100111101",
    954  => "010110010",
    955  => "001110011",
    956  => "111001101",
    957  => "001001100",
    958  => "011110101",
    959  => "011111011",
    960  => "000000111",
    961  => "010110101",
    962  => "000100001",
    963  => "100110000",
    964  => "111001101",
    965  => "111010110",
    966  => "000110100",
    967  => "001100001",
    968  => "011011001",
    969  => "010001100",
    970  => "100001100",
    971  => "100111000",
    972  => "101110100",
    973  => "011000111",
    974  => "010101101",
    975  => "101000100",
    976  => "011111101",
    977  => "011111100",
    978  => "110110101",
    979  => "000101010",
    980  => "110100101",
    981  => "011000101",
    982  => "011101101",
    983  => "100111110",
    984  => "111110001",
    985  => "011001001",
    986  => "101100110",
    987  => "100101011",
    988  => "110111111",
    989  => "101111001",
    990  => "001110011",
    991  => "101100010",
    992  => "000101101",
    993  => "001001011",
    994  => "100011001",
    995  => "011101001",
    996  => "010011010",
    997  => "011100111",
    998  => "100001110",
    999  => "110110011",
    1000 => "011101000",
    1001 => "000011101",
    1002 => "101100010",
    1003 => "111101001",
    1004 => "110110101",
    1005 => "101111011",
    1006 => "000100101",
    1007 => "010000011",
    1008 => "010010010",
    1009 => "110111110",
    1010 => "101101001",
    1011 => "011010111",
    1012 => "011111000",
    1013 => "011101111",
    1014 => "111010100",
    1015 => "010000000",
    1016 => "110111011",
    1017 => "110011110",
    1018 => "010001000",
    1019 => "000010101",
    1020 => "000111111",
    1021 => "111111010",
    1022 => "011111001",
    1023 => "011000011"
  );

  constant init_calendar_mem_512 : calendar_mem_type := (
    0   => "00000000000",
    1   => "11111111111",
    2   => "11111111111",
    3   => "11111111111",
    4   => "11111111111",
    5   => "11111111111",
    6   => "11111111111",
    7   => "11111111111",
    8   => "11111111111",
    9   => "11111111111",
    10  => "11111111111",
    11  => "11111111111",
    12  => "11111111111",
    13  => "11111111111",
    14  => "11111111111",
    15  => "11111111111",
    16  => "11111111111",
    17  => "11111111111",
    18  => "11111111111",
    19  => "11111111111",
    20  => "11111111111",
    21  => "11111111111",
    22  => "11111111111",
    23  => "11111111111",
    24  => "11111111111",
    25  => "11111111111",
    26  => "11111111111",
    27  => "11111111111",
    28  => "11111111111",
    29  => "11111111111",
    30  => "11111111111",
    31  => "11111111111",
    32  => "11111111111",
    33  => "11111111111",
    34  => "11111111111",
    35  => "11111111111",
    36  => "11111111111",
    37  => "11111111111",
    38  => "11111111111",
    39  => "11111111111",
    40  => "11111111111",
    41  => "11111111111",
    42  => "11111111111",
    43  => "11111111111",
    44  => "11111111111",
    45  => "11111111111",
    46  => "11111111111",
    47  => "11111111111",
    48  => "11111111111",
    49  => "11111111111",
    50  => "11111111111",
    51  => "11111111111",
    52  => "11111111111",
    53  => "11111111111",
    54  => "11111111111",
    55  => "11111111111",
    56  => "11111111111",
    57  => "11111111111",
    58  => "11111111111",
    59  => "11111111111",
    60  => "11111111111",
    61  => "11111111111",
    62  => "11111111111",
    63  => "11111111111",
    64  => "11111111111",
    65  => "11111111111",
    66  => "11111111111",
    67  => "11111111111",
    68  => "11111111111",
    69  => "11111111111",
    70  => "11111111111",
    71  => "11111111111",
    72  => "11111111111",
    73  => "11111111111",
    74  => "11111111111",
    75  => "11111111111",
    76  => "11111111111",
    77  => "11111111111",
    78  => "11111111111",
    79  => "11111111111",
    80  => "11111111111",
    81  => "11111111111",
    82  => "11111111111",
    83  => "11111111111",
    84  => "11111111111",
    85  => "11111111111",
    86  => "11111111111",
    87  => "11111111111",
    88  => "11111111111",
    89  => "11111111111",
    90  => "11111111111",
    91  => "11111111111",
    92  => "11111111111",
    93  => "11111111111",
    94  => "11111111111",
    95  => "11111111111",
    96  => "11111111111",
    97  => "11111111111",
    98  => "11111111111",
    99  => "11111111111",
    100 => "11111111111",
    101 => "11111111111",
    102 => "11111111111",
    103 => "11111111111",
    104 => "11111111111",
    105 => "11111111111",
    106 => "11111111111",
    107 => "11111111111",
    108 => "11111111111",
    109 => "11111111111",
    110 => "11111111111",
    111 => "11111111111",
    112 => "11111111111",
    113 => "11111111111",
    114 => "11111111111",
    115 => "11111111111",
    116 => "11111111111",
    117 => "11111111111",
    118 => "11111111111",
    119 => "11111111111",
    120 => "11111111111",
    121 => "11111111111",
    122 => "11111111111",
    123 => "11111111111",
    124 => "11111111111",
    125 => "11111111111",
    126 => "11111111111",
    127 => "11111111111",
    128 => "11111111111",
    129 => "11111111111",
    130 => "11111111111",
    131 => "11111111111",
    132 => "11111111111",
    133 => "11111111111",
    134 => "11111111111",
    135 => "11111111111",
    136 => "11111111111",
    137 => "11111111111",
    138 => "11111111111",
    139 => "11111111111",
    140 => "11111111111",
    141 => "11111111111",
    142 => "11111111111",
    143 => "11111111111",
    144 => "11111111111",
    145 => "11111111111",
    146 => "11111111111",
    147 => "11111111111",
    148 => "11111111111",
    149 => "11111111111",
    150 => "11111111111",
    151 => "11111111111",
    152 => "11111111111",
    153 => "11111111111",
    154 => "11111111111",
    155 => "11111111111",
    156 => "11111111111",
    157 => "11111111111",
    158 => "11111111111",
    159 => "11111111111",
    160 => "11111111111",
    161 => "11111111111",
    162 => "11111111111",
    163 => "11111111111",
    164 => "11111111111",
    165 => "11111111111",
    166 => "11111111111",
    167 => "11111111111",
    168 => "11111111111",
    169 => "11111111111",
    170 => "11111111111",
    171 => "11111111111",
    172 => "11111111111",
    173 => "11111111111",
    174 => "11111111111",
    175 => "11111111111",
    176 => "11111111111",
    177 => "11111111111",
    178 => "11111111111",
    179 => "11111111111",
    180 => "11111111111",
    181 => "11111111111",
    182 => "11111111111",
    183 => "11111111111",
    184 => "11111111111",
    185 => "11111111111",
    186 => "11111111111",
    187 => "11111111111",
    188 => "11111111111",
    189 => "11111111111",
    190 => "11111111111",
    191 => "11111111111",
    192 => "11111111111",
    193 => "11111111111",
    194 => "11111111111",
    195 => "11111111111",
    196 => "11111111111",
    197 => "11111111111",
    198 => "11111111111",
    199 => "11111111111",
    200 => "11111111111",
    201 => "11111111111",
    202 => "11111111111",
    203 => "11111111111",
    204 => "11111111111",
    205 => "11111111111",
    206 => "11111111111",
    207 => "11111111111",
    208 => "11111111111",
    209 => "11111111111",
    210 => "11111111111",
    211 => "11111111111",
    212 => "11111111111",
    213 => "11111111111",
    214 => "11111111111",
    215 => "11111111111",
    216 => "11111111111",
    217 => "11111111111",
    218 => "11111111111",
    219 => "11111111111",
    220 => "11111111111",
    221 => "11111111111",
    222 => "11111111111",
    223 => "11111111111",
    224 => "11111111111",
    225 => "11111111111",
    226 => "11111111111",
    227 => "11111111111",
    228 => "11111111111",
    229 => "11111111111",
    230 => "11111111111",
    231 => "11111111111",
    232 => "11111111111",
    233 => "11111111111",
    234 => "11111111111",
    235 => "11111111111",
    236 => "11111111111",
    237 => "11111111111",
    238 => "11111111111",
    239 => "11111111111",
    240 => "11111111111",
    241 => "11111111111",
    242 => "11111111111",
    243 => "11111111111",
    244 => "11111111111",
    245 => "11111111111",
    246 => "11111111111",
    247 => "11111111111",
    248 => "11111111111",
    249 => "11111111111",
    250 => "11111111111",
    251 => "11111111111",
    252 => "11111111111",
    253 => "11111111111",
    254 => "11111111111",
    255 => "11111111111",
    256 => "11111111111",
    257 => "11111111111",
    258 => "11111111111",
    259 => "11111111111",
    260 => "11111111111",
    261 => "11111111111",
    262 => "11111111111",
    263 => "11111111111",
    264 => "11111111111",
    265 => "11111111111",
    266 => "11111111111",
    267 => "11111111111",
    268 => "11111111111",
    269 => "11111111111",
    270 => "11111111111",
    271 => "11111111111",
    272 => "11111111111",
    273 => "11111111111",
    274 => "11111111111",
    275 => "11111111111",
    276 => "11111111111",
    277 => "11111111111",
    278 => "11111111111",
    279 => "11111111111",
    280 => "11111111111",
    281 => "11111111111",
    282 => "11111111111",
    283 => "11111111111",
    284 => "11111111111",
    285 => "11111111111",
    286 => "11111111111",
    287 => "11111111111",
    288 => "11111111111",
    289 => "11111111111",
    290 => "11111111111",
    291 => "11111111111",
    292 => "11111111111",
    293 => "11111111111",
    294 => "11111111111",
    295 => "11111111111",
    296 => "11111111111",
    297 => "11111111111",
    298 => "11111111111",
    299 => "11111111111",
    300 => "11111111111",
    301 => "11111111111",
    302 => "11111111111",
    303 => "11111111111",
    304 => "11111111111",
    305 => "11111111111",
    306 => "11111111111",
    307 => "11111111111",
    308 => "11111111111",
    309 => "11111111111",
    310 => "11111111111",
    311 => "11111111111",
    312 => "11111111111",
    313 => "11111111111",
    314 => "11111111111",
    315 => "11111111111",
    316 => "11111111111",
    317 => "11111111111",
    318 => "11111111111",
    319 => "11111111111",
    320 => "11111111111",
    321 => "11111111111",
    322 => "11111111111",
    323 => "11111111111",
    324 => "11111111111",
    325 => "11111111111",
    326 => "11111111111",
    327 => "11111111111",
    328 => "11111111111",
    329 => "11111111111",
    330 => "11111111111",
    331 => "11111111111",
    332 => "11111111111",
    333 => "11111111111",
    334 => "11111111111",
    335 => "11111111111",
    336 => "11111111111",
    337 => "11111111111",
    338 => "11111111111",
    339 => "11111111111",
    340 => "11111111111",
    341 => "11111111111",
    342 => "11111111111",
    343 => "11111111111",
    344 => "11111111111",
    345 => "11111111111",
    346 => "11111111111",
    347 => "11111111111",
    348 => "11111111111",
    349 => "11111111111",
    350 => "11111111111",
    351 => "11111111111",
    352 => "11111111111",
    353 => "11111111111",
    354 => "11111111111",
    355 => "11111111111",
    356 => "11111111111",
    357 => "11111111111",
    358 => "11111111111",
    359 => "11111111111",
    360 => "11111111111",
    361 => "11111111111",
    362 => "11111111111",
    363 => "11111111111",
    364 => "11111111111",
    365 => "11111111111",
    366 => "11111111111",
    367 => "11111111111",
    368 => "11111111111",
    369 => "11111111111",
    370 => "11111111111",
    371 => "11111111111",
    372 => "11111111111",
    373 => "11111111111",
    374 => "11111111111",
    375 => "11111111111",
    376 => "11111111111",
    377 => "11111111111",
    378 => "11111111111",
    379 => "11111111111",
    380 => "11111111111",
    381 => "11111111111",
    382 => "11111111111",
    383 => "11111111111",
    384 => "11111111111",
    385 => "11111111111",
    386 => "11111111111",
    387 => "11111111111",
    388 => "11111111111",
    389 => "11111111111",
    390 => "11111111111",
    391 => "11111111111",
    392 => "11111111111",
    393 => "11111111111",
    394 => "11111111111",
    395 => "11111111111",
    396 => "11111111111",
    397 => "11111111111",
    398 => "11111111111",
    399 => "11111111111",
    400 => "11111111111",
    401 => "11111111111",
    402 => "11111111111",
    403 => "11111111111",
    404 => "11111111111",
    405 => "11111111111",
    406 => "11111111111",
    407 => "11111111111",
    408 => "11111111111",
    409 => "11111111111",
    410 => "11111111111",
    411 => "11111111111",
    412 => "11111111111",
    413 => "11111111111",
    414 => "11111111111",
    415 => "11111111111",
    416 => "11111111111",
    417 => "11111111111",
    418 => "11111111111",
    419 => "11111111111",
    420 => "11111111111",
    421 => "11111111111",
    422 => "11111111111",
    423 => "11111111111",
    424 => "11111111111",
    425 => "11111111111",
    426 => "11111111111",
    427 => "11111111111",
    428 => "11111111111",
    429 => "11111111111",
    430 => "11111111111",
    431 => "11111111111",
    432 => "11111111111",
    433 => "11111111111",
    434 => "11111111111",
    435 => "11111111111",
    436 => "11111111111",
    437 => "11111111111",
    438 => "11111111111",
    439 => "11111111111",
    440 => "11111111111",
    441 => "11111111111",
    442 => "11111111111",
    443 => "11111111111",
    444 => "11111111111",
    445 => "11111111111",
    446 => "11111111111",
    447 => "11111111111",
    448 => "11111111111",
    449 => "11111111111",
    450 => "11111111111",
    451 => "11111111111",
    452 => "11111111111",
    453 => "11111111111",
    454 => "11111111111",
    455 => "11111111111",
    456 => "11111111111",
    457 => "11111111111",
    458 => "11111111111",
    459 => "11111111111",
    460 => "11111111111",
    461 => "11111111111",
    462 => "11111111111",
    463 => "11111111111",
    464 => "11111111111",
    465 => "11111111111",
    466 => "11111111111",
    467 => "11111111111",
    468 => "11111111111",
    469 => "11111111111",
    470 => "11111111111",
    471 => "11111111111",
    472 => "11111111111",
    473 => "11111111111",
    474 => "11111111111",
    475 => "11111111111",
    476 => "11111111111",
    477 => "11111111111",
    478 => "11111111111",
    479 => "11111111111",
    480 => "11111111111",
    481 => "11111111111",
    482 => "11111111111",
    483 => "11111111111",
    484 => "11111111111",
    485 => "11111111111",
    486 => "11111111111",
    487 => "11111111111",
    488 => "11111111111",
    489 => "11111111111",
    490 => "11111111111",
    491 => "11111111111",
    492 => "11111111111",
    493 => "11111111111",
    494 => "11111111111",
    495 => "11111111111",
    496 => "11111111111",
    497 => "11111111111",
    498 => "11111111111",
    499 => "11111111111",
    500 => "11111111111",
    501 => "11111111111",
    502 => "11111111111",
    503 => "11111111111",
    504 => "11111111111",
    505 => "11111111111",
    506 => "11111111111",
    507 => "11111111111",
    508 => "11111111111",
    509 => "11111111111",
    510 => "11111111111",
    511 => "11111111111"
  );

end package;
