-- RP simulation package
library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use ieee.numeric_std.all;
  use work.constants_pkg.all; -- Import constants

package bram_init_pkg is

  -- Memory
  type rate_mem_type is array (0 to 2 ** 6 - 1) of std_logic_vector(16 - 1 downto 0);
  type RP_mem_type is array (0 to 2 ** 6 - 1) of std_logic_vector(105 - 1 downto 0);

  constant init_rate_mem_16 : rate_mem_type := (
    0  => "0000000000000111", -- 7
    1  => "0000000000000111", -- 7
    2  => "0000000000000111", -- 7
    3  => "0000000000000111", -- 7
    4  => "0000000000000111", -- 7
    5  => "0000000000000111", -- 7
    6  => "0000000000000111", -- 7
    7  => "0000000000000111", -- 7
    8  => "0000000000000111", -- 7
    9  => "0000000000000110", -- 6
    10 => "0000000000000110", -- 6
    11 => "0000000000000110", -- 6
    12 => "0000000000000111", -- 7
    13 => "0000000000000111", -- 7
    14 => "0000000000000111", -- 7
    15 => "0000000000000111", -- 7
    16 => "0000000000000111", -- 7
    17 => "0000000000000111", -- 7
    18 => "0000000000000111", -- 7
    19 => "0000000000000111", -- 7
    20 => "0000000000000111", -- 7
    21 => "0000000000000111", -- 7
    22 => "0000000000000111", -- 7
    23 => "0000000000000111", -- 7
    24 => "0000000000000111", -- 7
    25 => "0000000000000111", -- 7
    26 => "0000000000000111", -- 7
    27 => "0000000000000111", -- 7
    28 => "0000000000000111", -- 7
    29 => "0000000000000111", -- 7
    30 => "0000000000000111", -- 7
    31 => "0000000000000111", -- 7
    32 => "0000000000000111", -- 7
    33 => "0000000000000111", -- 7
    34 => "0000000000000111", -- 7
    35 => "0000000000000111", -- 7
    36 => "0000000000000111", -- 7
    37 => "0000000000000111", -- 7
    38 => "0000000000000111", -- 7
    39 => "0000000000000111", -- 7
    40 => "0000000000000111", -- 7
    41 => "0000000000000111", -- 7
    42 => "0000000000000111", -- 7
    43 => "0000000000000111", -- 7
    44 => "0000000000000111", -- 7
    45 => "0000000000000111", -- 7
    46 => "0000000000000111", -- 7
    47 => "0000000000000111", -- 7
    48 => "0000000000000111", -- 7
    49 => "0000000000000111", -- 7
    50 => "0000000000000111", -- 7
    51 => "0000000000000111", -- 7
    52 => "0000000000000111", -- 7
    53 => "0000000000000111", -- 7
    54 => "0000000000000111", -- 7
    55 => "0000000000000111", -- 7
    56 => "0000000000000111", -- 7
    57 => "0000000000000111", -- 7
    58 => "0000000000000111", -- 7
    59 => "0000000000000111", -- 7
    60 => "0000000000000111", -- 7
    61 => "0000000000000111", -- 7
    62 => "0000000000000111", -- 7
    63 => "0000000000000111" -- 7
  );

  constant init_RP_mem_16 : RP_mem_type := (
    0  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    1  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    2  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    3  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    4  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    5  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    6  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    7  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    8  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    9  => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    10 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    11 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    12 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    13 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    14 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    15 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    16 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    17 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    18 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    19 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    20 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    21 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    22 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    23 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    24 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    25 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    26 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    27 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    28 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    29 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    30 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    31 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    32 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    33 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    34 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    35 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    36 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    37 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    38 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    39 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    40 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    41 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    42 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    43 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    44 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    45 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    46 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    47 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    48 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    49 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    50 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    51 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    52 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    53 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    54 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    55 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    56 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    57 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    58 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    59 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    60 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    61 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    62 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111",
    63 => "000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110111111111111111"
  );

end package;
