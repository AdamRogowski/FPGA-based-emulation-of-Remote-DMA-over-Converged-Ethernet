library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use ieee.numeric_std.all;
  use work.constants_pkg.all;

package flow_array_pkg is

  type FlowEntry is record
    flow_addr : std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0);
    max_rate  : unsigned(RATE_BIT_RESOLUTION_WIDTH - 1 downto 0);
    cur_rate  : unsigned(RATE_BIT_RESOLUTION_WIDTH - 1 downto 0);
  end record;

  type FlowArray is array (0 to NUM_FLOWS_TOTAL - 1) of FlowEntry;

  -- When changing the flow array, update constants_pkg.vhd to match the new flow array size
  -- Update:
  -- NUM_GROUPS
  -- NUM_FLOWS
  -- FLAT_FLOW_ADDRESS_WIDTH

  -- If rate resolution is changed, update the following constants in constants_pkg.vhd:
  -- RATE_BIT_RESOLUTION
  -- RATE_BIT_RESOLUTION_WIDTH
  constant FLOWS : FlowArray := (
    0   => ("000000000", "1111111111", "0110111100"),
    1   => ("000000001", "1111111111", "1010010000"),
    2   => ("000000010", "1111111111", "0000010010"),
    3   => ("000000011", "1111111111", "1101101011"),
    4   => ("000000100", "1111111111", "1010110001"),
    5   => ("000000101", "1111111111", "1100100011"),
    6   => ("000000110", "1111111111", "0010001000"),
    7   => ("000000111", "1111111111", "1100110110"),
    8   => ("000001000", "1111111111", "1100101111"),
    9   => ("000001001", "1111111111", "0110001101"),
    10  => ("000001010", "1111111111", "0000110000"),
    11  => ("000001011", "1111111111", "1101001100"),
    12  => ("000001100", "1111111111", "1110000111"),
    13  => ("000001101", "1111111111", "1110001011"),
    14  => ("000001110", "1111111111", "1111101110"),
    15  => ("000001111", "1111111111", "0101100111"),
    16  => ("000010000", "1111111111", "1001011101"),
    17  => ("000010001", "1111111111", "0010110110"),
    18  => ("000010010", "1111111111", "0111001010"),
    19  => ("000010011", "1111111111", "1001011011"),
    20  => ("000010100", "1111111111", "1111111001"),
    21  => ("000010101", "1111111111", "0001101100"),
    22  => ("000010110", "1111111111", "0110111011"),
    23  => ("000010111", "1111111111", "1001001110"),
    24  => ("000011000", "1111111111", "0101111101"),
    25  => ("000011001", "1111111111", "0111010111"),
    26  => ("000011010", "1111111111", "0000100110"),
    27  => ("000011011", "1111111111", "1100111011"),
    28  => ("000011100", "1111111111", "1000000100"),
    29  => ("000011101", "1111111111", "1010011101"),
    30  => ("000011110", "1111111111", "1001001101"),
    31  => ("000011111", "1111111111", "0001110011"),
    32  => ("000100000", "1111111111", "0010010000"),
    33  => ("000100001", "1111111111", "0000110011"),
    34  => ("000100010", "1111111111", "1010101101"),
    35  => ("000100011", "1111111111", "0101111000"),
    36  => ("000100100", "1111111111", "0110010011"),
    37  => ("000100101", "1111111111", "1110100010"),
    38  => ("000100110", "1111111111", "1110110101"),
    39  => ("000100111", "1111111111", "1010011010"),
    40  => ("000101000", "1111111111", "1001000010"),
    41  => ("000101001", "1111111111", "1100111100"),
    42  => ("000101010", "1111111111", "1001111011"),
    43  => ("000101011", "1111111111", "0000101111"),
    44  => ("000101100", "1111111111", "1000110000"),
    45  => ("000101101", "1111111111", "0101100100"),
    46  => ("000101110", "1111111111", "1111100100"),
    47  => ("000101111", "1111111111", "1110110100"),
    48  => ("000110000", "1111111111", "1001111000"),
    49  => ("000110001", "1111111111", "0000101001"),
    50  => ("000110010", "1111111111", "0111101111"),
    51  => ("000110011", "1111111111", "1011110001"),
    52  => ("000110100", "1111111111", "1010101101"),
    53  => ("000110101", "1111111111", "1101011101"),
    54  => ("000110110", "1111111111", "0111011000"),
    55  => ("000110111", "1111111111", "1000011001"),
    56  => ("000111000", "1111111111", "0111100100"),
    57  => ("000111001", "1111111111", "0100010010"),
    58  => ("000111010", "1111111111", "1010101001"),
    59  => ("000111011", "1111111111", "1101101110"),
    60  => ("000111100", "1111111111", "0100110010"),
    61  => ("000111101", "1111111111", "0110010010"),
    62  => ("000111110", "1111111111", "1100100010"),
    63  => ("000111111", "1111111111", "1010011111"),
    64  => ("001000000", "1111111111", "0000001001"),
    65  => ("001000001", "1111111111", "0100000111"),
    66  => ("001000010", "1111111111", "1001000111"),
    67  => ("001000011", "1111111111", "0011000010"),
    68  => ("001000100", "1111111111", "1110110100"),
    69  => ("001000101", "1111111111", "1000010010"),
    70  => ("001000110", "1111111111", "0010000011"),
    71  => ("001000111", "1111111111", "1101001101"),
    72  => ("001001000", "1111111111", "1000111111"),
    73  => ("001001001", "1111111111", "1101010011"),
    74  => ("001001010", "1111111111", "0000010100"),
    75  => ("001001011", "1111111111", "0011101011"),
    76  => ("001001100", "1111111111", "1000011010"),
    77  => ("001001101", "1111111111", "0011000010"),
    78  => ("001001110", "1111111111", "1010110010"),
    79  => ("001001111", "1111111111", "0101011110"),
    80  => ("001010000", "1111111111", "1011111110"),
    81  => ("001010001", "1111111111", "1010011101"),
    82  => ("001010010", "1111111111", "0100110100"),
    83  => ("001010011", "1111111111", "1100111110"),
    84  => ("001010100", "1111111111", "0010010001"),
    85  => ("001010101", "1111111111", "1001000010"),
    86  => ("001010110", "1111111111", "0001100111"),
    87  => ("001010111", "1111111111", "0011001011"),
    88  => ("001011000", "1111111111", "1011101010"),
    89  => ("001011001", "1111111111", "1000011110"),
    90  => ("001011010", "1111111111", "1000101110"),
    91  => ("001011011", "1111111111", "1100110111"),
    92  => ("001011100", "1111111111", "1000111011"),
    93  => ("001011101", "1111111111", "0011111000"),
    94  => ("001011110", "1111111111", "1000000100"),
    95  => ("001011111", "1111111111", "0011000101"),
    96  => ("001100000", "1111111111", "1000100110"),
    97  => ("001100001", "1111111111", "1101001110"),
    98  => ("001100010", "1111111111", "1110010110"),
    99  => ("001100011", "1111111111", "0001110110"),
    100 => ("001100100", "1111111111", "1000001011"),
    101 => ("001100101", "1111111111", "0111010010"),
    102 => ("001100110", "1111111111", "1001011001"),
    103 => ("001100111", "1111111111", "1011011000"),
    104 => ("001101000", "1111111111", "0011001010"),
    105 => ("001101001", "1111111111", "0011010001"),
    106 => ("001101010", "1111111111", "1010110110"),
    107 => ("001101011", "1111111111", "1001100010"),
    108 => ("001101100", "1111111111", "0100101111"),
    109 => ("001101101", "1111111111", "0011001000"),
    110 => ("001101110", "1111111111", "0001001011"),
    111 => ("001101111", "1111111111", "0000100100"),
    112 => ("001110000", "1111111111", "0000100000"),
    113 => ("001110001", "1111111111", "1011001100"),
    114 => ("001110010", "1111111111", "0100000010"),
    115 => ("001110011", "1111111111", "1100001110"),
    116 => ("001110100", "1111111111", "0101111100"),
    117 => ("001110101", "1111111111", "1011010001"),
    118 => ("001110110", "1111111111", "0111111001"),
    119 => ("001110111", "1111111111", "0111110011"),
    120 => ("001111000", "1111111111", "0001000010"),
    121 => ("001111001", "1111111111", "1110000110"),
    122 => ("001111010", "1111111111", "1001001010"),
    123 => ("001111011", "1111111111", "1100111100"),
    124 => ("001111100", "1111111111", "0001001101"),
    125 => ("001111101", "1111111111", "0011110110"),
    126 => ("001111110", "1111111111", "0100011010"),
    127 => ("001111111", "1111111111", "1001110000"),
    128 => ("010000000", "1111111111", "1001001011"),
    129 => ("010000001", "1111111111", "0110011001"),
    130 => ("010000010", "1111111111", "1110001111"),
    131 => ("010000011", "1111111111", "0001010101"),
    132 => ("010000100", "1111111111", "0011101101"),
    133 => ("010000101", "1111111111", "1011100111"),
    134 => ("010000110", "1111111111", "1000100110"),
    135 => ("010000111", "1111111111", "1110011100"),
    136 => ("010001000", "1111111111", "0010110011"),
    137 => ("010001001", "1111111111", "1001011011"),
    138 => ("010001010", "1111111111", "0111110000"),
    139 => ("010001011", "1111111111", "1100111001"),
    140 => ("010001100", "1111111111", "0000111000"),
    141 => ("010001101", "1111111111", "0011101111"),
    142 => ("010001110", "1111111111", "0011000001"),
    143 => ("010001111", "1111111111", "1100110111"),
    144 => ("010010000", "1111111111", "1001111011"),
    145 => ("010010001", "1111111111", "1010011010"),
    146 => ("010010010", "1111111111", "0010101100"),
    147 => ("010010011", "1111111111", "1010001010"),
    148 => ("010010100", "1111111111", "0110011110"),
    149 => ("010010101", "1111111111", "1100110111"),
    150 => ("010010110", "1111111111", "0110111110"),
    151 => ("010010111", "1111111111", "1010110111"),
    152 => ("010011000", "1111111111", "1010001011"),
    153 => ("010011001", "1111111111", "1000000100"),
    154 => ("010011010", "1111111111", "1010010111"),
    155 => ("010011011", "1111111111", "1001111001"),
    156 => ("010011100", "1111111111", "0010101111"),
    157 => ("010011101", "1111111111", "0010111111"),
    158 => ("010011110", "1111111111", "0111101111"),
    159 => ("010011111", "1111111111", "1000111011"),
    160 => ("010100000", "1111111111", "0001000100"),
    161 => ("010100001", "1111111111", "0001110101"),
    162 => ("010100010", "1111111111", "1111010001"),
    163 => ("010100011", "1111111111", "0101011001"),
    164 => ("010100100", "1111111111", "0101101111"),
    165 => ("010100101", "1111111111", "1100100000"),
    166 => ("010100110", "1111111111", "0100001111"),
    167 => ("010100111", "1111111111", "0101111100"),
    168 => ("010101000", "1111111111", "0010100100"),
    169 => ("010101001", "1111111111", "1000011010"),
    170 => ("010101010", "1111111111", "1011110101"),
    171 => ("010101011", "1111111111", "1001000000"),
    172 => ("010101100", "1111111111", "0001011010"),
    173 => ("010101101", "1111111111", "1010011011"),
    174 => ("010101110", "1111111111", "1001000011"),
    175 => ("010101111", "1111111111", "1000101101"),
    176 => ("010110000", "1111111111", "0001101010"),
    177 => ("010110001", "1111111111", "0011101101"),
    178 => ("010110010", "1111111111", "1000000110"),
    179 => ("010110011", "1111111111", "1001100111"),
    180 => ("010110100", "1111111111", "1110011011"),
    181 => ("010110101", "1111111111", "1001000101"),
    182 => ("010110110", "1111111111", "0000011100"),
    183 => ("010110111", "1111111111", "1001110111"),
    184 => ("010111000", "1111111111", "0111011100"),
    185 => ("010111001", "1111111111", "0000011000"),
    186 => ("010111010", "1111111111", "0000010010"),
    187 => ("010111011", "1111111111", "0100111010"),
    188 => ("010111100", "1111111111", "0101001011"),
    189 => ("010111101", "1111111111", "0011101110"),
    190 => ("010111110", "1111111111", "0100000011"),
    191 => ("010111111", "1111111111", "1101011001"),
    192 => ("011000000", "1111111111", "1100001011"),
    193 => ("011000001", "1111111111", "1001101111"),
    194 => ("011000010", "1111111111", "1100100100"),
    195 => ("011000011", "1111111111", "0010011000"),
    196 => ("011000100", "1111111111", "0001100110"),
    197 => ("011000101", "1111111111", "1010100100"),
    198 => ("011000110", "1111111111", "0010110010"),
    199 => ("011000111", "1111111111", "1111010110"),
    200 => ("011001000", "1111111111", "1101111101"),
    201 => ("011001001", "1111111111", "0010010011"),
    202 => ("011001010", "1111111111", "0110101000"),
    203 => ("011001011", "1111111111", "0101101001"),
    204 => ("011001100", "1111111111", "0100000011"),
    205 => ("011001101", "1111111111", "1000001011"),
    206 => ("011001110", "1111111111", "0001010001"),
    207 => ("011001111", "1111111111", "1111100110"),
    208 => ("011010000", "1111111111", "0011010001"),
    209 => ("011010001", "1111111111", "0001101010"),
    210 => ("011010010", "1111111111", "1110110111"),
    211 => ("011010011", "1111111111", "0100111111"),
    212 => ("011010100", "1111111111", "1100010011"),
    213 => ("011010101", "1111111111", "1000000110"),
    214 => ("011010110", "1111111111", "0000011111"),
    215 => ("011010111", "1111111111", "1110111111"),
    216 => ("011011000", "1111111111", "0000100110"),
    217 => ("011011001", "1111111111", "0011000100"),
    218 => ("011011010", "1111111111", "1011100111"),
    219 => ("011011011", "1111111111", "0110101001"),
    220 => ("011011100", "1111111111", "1010011000"),
    221 => ("011011101", "1111111111", "0101001101"),
    222 => ("011011110", "1111111111", "1110101111"),
    223 => ("011011111", "1111111111", "0010111000"),
    224 => ("011100000", "1111111111", "1000110111"),
    225 => ("011100001", "1111111111", "0110001110"),
    226 => ("011100010", "1111111111", "0101100000"),
    227 => ("011100011", "1111111111", "1111001000"),
    228 => ("011100100", "1111111111", "0101011000"),
    229 => ("011100101", "1111111111", "1100001011"),
    230 => ("011100110", "1111111111", "1010011000"),
    231 => ("011100111", "1111111111", "0011100100"),
    232 => ("011101000", "1111111111", "1010000110"),
    233 => ("011101001", "1111111111", "0011111011"),
    234 => ("011101010", "1111111111", "1110010100"),
    235 => ("011101011", "1111111111", "0001111100"),
    236 => ("011101100", "1111111111", "0010100001"),
    237 => ("011101101", "1111111111", "1111000010"),
    238 => ("011101110", "1111111111", "0011000000"),
    239 => ("011101111", "1111111111", "0101110011"),
    240 => ("011110000", "1111111111", "0111100011"),
    241 => ("011110001", "1111111111", "0100001000"),
    242 => ("011110010", "1111111111", "0011110000"),
    243 => ("011110011", "1111111111", "0100111111"),
    244 => ("011110100", "1111111111", "1111010011"),
    245 => ("011110101", "1111111111", "1101110010"),
    246 => ("011110110", "1111111111", "0010000011"),
    247 => ("011110111", "1111111111", "0101101100"),
    248 => ("011111000", "1111111111", "1111001011"),
    249 => ("011111001", "1111111111", "0010110101"),
    250 => ("011111010", "1111111111", "1000111101"),
    251 => ("011111011", "1111111111", "0000000100"),
    252 => ("011111100", "1111111111", "1111100100"),
    253 => ("011111101", "1111111111", "0110101011"),
    254 => ("011111110", "1111111111", "0101111011"),
    255 => ("011111111", "1111111111", "1011101111")
  );

end package;
