-- divider.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
library divider_lpm_divide_201;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity divider is
	port (
		numer    : in  std_logic_vector(35 downto 0) := (others => '0'); --  lpm_divide_input.numer
		denom    : in  std_logic_vector(15 downto 0) := (others => '0'); --                  .denom
		clock    : in  std_logic                     := '0';             --                  .clock
		quotient : out std_logic_vector(35 downto 0);                    -- lpm_divide_output.quotient
		remain   : out std_logic_vector(15 downto 0)                     --                  .remain
	);
end entity divider;

architecture rtl of divider is
	component divider_lpm_divide_201_gohehnq is
		port (
			numer    : in  std_logic_vector(35 downto 0) := (others => 'X'); -- numer
			denom    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- denom
			clock    : in  std_logic                     := 'X';             -- clock
			quotient : out std_logic_vector(35 downto 0);                    -- quotient
			remain   : out std_logic_vector(15 downto 0)                     -- remain
		);
	end component divider_lpm_divide_201_gohehnq;

	for lpm_divide_0 : divider_lpm_divide_201_gohehnq
		use entity divider_lpm_divide_201.divider_lpm_divide_201_gohehnq;
begin

	lpm_divide_0 : component divider_lpm_divide_201_gohehnq
		port map (
			numer    => numer,    --  lpm_divide_input.numer
			denom    => denom,    --                  .denom
			clock    => clock,    --                  .clock
			quotient => quotient, -- lpm_divide_output.quotient
			remain   => remain    --                  .remain
		);

end architecture rtl; -- of divider
