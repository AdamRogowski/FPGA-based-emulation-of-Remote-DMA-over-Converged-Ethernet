-- RP simulation package
library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use ieee.numeric_std.all;
  use work.constants_pkg.all; -- Import constants

package bram_init_pkg is

  -- Memory
  type rate_mem_type is array (0 to 2 ** 6 - 1) of std_logic_vector(17 - 1 downto 0);
  type RP_mem_type is array (0 to 2 ** 6 - 1) of std_logic_vector(111 - 1 downto 0);

  constant init_rate_mem_16 : rate_mem_type := (
    0  => "00010110010111001", -- 7 
    1  => "00010110010111001", -- 7
    2  => "00010110010111001", -- 7
    3  => "00010110010111001", -- 7
    4  => "00010110010111001", -- 7
    5  => "00010110010111001", -- 7
    6  => "00010110010111001", -- 7
    7  => "00010110010111001", -- 7
    8  => "00010110010111001", -- 7
    9  => "00010110010111001", -- 6
    10 => "00010110010111001", -- 6
    11 => "00010110010111001", -- 6
    12 => "00010110010111001", -- 7
    13 => "00010110010111001", -- 7
    14 => "00010110010111001", -- 7
    15 => "00010110010111001", -- 7
    16 => "00010110010111001", -- 7
    17 => "00010110010111001", -- 7
    18 => "00010110010111001", -- 7
    19 => "00010110010111001", -- 7
    20 => "00010110010111001", -- 7
    21 => "00010110010111001", -- 7
    22 => "00010110010111001", -- 7
    23 => "00010110010111001", -- 7
    24 => "00010110010111001", -- 7
    25 => "00010110010111001", -- 7
    26 => "00010110010111001", -- 7
    27 => "00010110010111001", -- 7
    28 => "00010110010111001", -- 7
    29 => "00010110010111001", -- 7
    30 => "00010110010111001", -- 7
    31 => "00010110010111001", -- 7
    32 => "00010110010111001", -- 7
    33 => "00010110010111001", -- 7
    34 => "00010110010111001", -- 7
    35 => "00010110010111001", -- 7
    36 => "00010110010111001", -- 7
    37 => "00010110010111001", -- 7
    38 => "00010110010111001", -- 7
    39 => "00010110010111001", -- 7
    40 => "00010110010111001", -- 7
    41 => "00010110010111001", -- 7
    42 => "00010110010111001", -- 7
    43 => "00010110010111001", -- 7
    44 => "00010110010111001", -- 7
    45 => "00010110010111001", -- 7
    46 => "00010110010111001", -- 7
    47 => "00010110010111001", -- 7
    48 => "00010110010111001", -- 7
    49 => "00010110010111001", -- 7
    50 => "00010110010111001", -- 7
    51 => "00010110010111001", -- 7
    52 => "00000000000001011", -- 7
    53 => "00010110010111001", -- 7
    54 => "00010110010111001", -- 7
    55 => "00010110010111001", -- 7
    56 => "00010110010111001", -- 7
    57 => "00010110010111001", -- 7
    58 => "00010110010111001", -- 7
    59 => "00010110010111001", -- 7
    60 => "00010110010111001", -- 7
    61 => "00010110010111001", -- 7
    62 => "00010110010111001", -- 7
    63 => "00010110010111001" -- 7
  );

  constant init_RP_mem_16 : RP_mem_type := (
    0  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000011111111111011111111111111111",
    1  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    2  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    3  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    4  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    5  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    6  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    7  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    8  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    9  => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    10 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    11 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    12 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    13 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    14 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    15 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    16 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    17 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    18 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    19 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    20 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    21 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    22 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    23 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    24 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    25 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    26 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    27 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    28 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    29 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    30 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    31 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    32 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    33 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    34 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    35 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    36 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    37 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    38 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    39 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    40 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    41 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    42 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    43 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    44 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    45 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    46 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    47 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    48 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    49 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    50 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    51 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    52 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    53 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    54 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    55 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    56 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    57 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    58 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    59 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    60 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    61 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    62 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111",
    63 => "000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111111011111111111111111"
  );

end package;
