library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use ieee.numeric_std.all;
  use work.constants_pkg.all;

package flow_array_pkg is

  type FlowEntry is record
    flow_addr : std_logic_vector(FLOW_ADDRESS_WIDTH - 1 downto 0);
    max_rate  : unsigned(RATE_BIT_RESOLUTION_WIDTH - 1 downto 0);
    cur_rate  : unsigned(RATE_BIT_RESOLUTION_WIDTH - 1 downto 0);
  end record;

  type FlowArray is array (0 to NUM_FLOWS_TOTAL - 1) of FlowEntry;

  -- When changing the flow array, update constants_pkg.vhd to match the new flow array size
  -- Update:
  -- NUM_GROUPS
  -- NUM_FLOWS
  -- FLAT_FLOW_ADDRESS_WIDTH

  -- If rate resolution is changed, update the following constants in constants_pkg.vhd:
  -- RATE_BIT_RESOLUTION
  -- RATE_BIT_RESOLUTION_WIDTH
  constant FLOWS : FlowArray := (
    0   => ("000000000", "00000000000001010", "11100010110110100"),
    1   => ("000000001", "00000000000001010", "00111111100101101"),
    2   => ("000000010", "00000000000001010", "01001101010011111"),
    3   => ("000000011", "00000000000001010", "10100110111100001"),
    4   => ("000000100", "00000000000001010", "01101011000111010"),
    5   => ("000000101", "00000000000001010", "01011100001110010"),
    6   => ("000000110", "00000000000001010", "11001101111011000"),
    7   => ("000000111", "00000000000001010", "01111001000110111"),
    8   => ("000001000", "00000000000001010", "00000111010000001"),
    9   => ("000001001", "00000000000001010", "10111101110101011"),
    10  => ("000001010", "00000000000001010", "01110000101101110"),
    11  => ("000001011", "00000000000001010", "01011111100010111"),
    12  => ("000001100", "00000000000001010", "11110100011000100"),
    13  => ("000001101", "00000000000001010", "00010101111111100"),
    14  => ("000001110", "00000000000001010", "01101010000000101"),
    15  => ("000001111", "00000000000001010", "00001100010110010"),
    16  => ("000010000", "00000000000001010", "10001000100101010"),
    17  => ("000010001", "00000000000001010", "01010011111011111"),
    18  => ("000010010", "00000000000001010", "10110001110001000"),
    19  => ("000010011", "00000000000001010", "01100110100001010"),
    20  => ("000010100", "00000000000001010", "10001000101001101"),
    21  => ("000010101", "00000000000001010", "10110101111011100"),
    22  => ("000010110", "00000000000001010", "01000011000111101"),
    23  => ("000010111", "00000000000001010", "01001011100011011"),
    24  => ("000011000", "00000000000001010", "00111011001110011"),
    25  => ("000011001", "00000000000001010", "01000001110011010"),
    26  => ("000011010", "00000000000001010", "00111001001100101"),
    27  => ("000011011", "00000000000001010", "11101001011011011"),
    28  => ("000011100", "00000000000001010", "11111001111100000"),
    29  => ("000011101", "00000000000001010", "00101100111111111"),
    30  => ("000011110", "00000000000001010", "10111111011010101"),
    31  => ("000011111", "00000000000001010", "01010010111001101"),
    32  => ("000100000", "00000000000001010", "10111010001011001"),
    33  => ("000100001", "00000000000001010", "11011010011101101"),
    34  => ("000100010", "00000000000001010", "11111011100000010"),
    35  => ("000100011", "00000000000001010", "00100001010101111"),
    36  => ("000100100", "00000000000001010", "10010100000001100"),
    37  => ("000100101", "00000000000001010", "10111101011001000"),
    38  => ("000100110", "00000000000001010", "00100100011011000"),
    39  => ("000100111", "00000000000001010", "11010111001111111"),
    40  => ("000101000", "00000000000001010", "11010111101011110"),
    41  => ("000101001", "00000000000001010", "00101000011100010"),
    42  => ("000101010", "00000000000001010", "00011000001110110"),
    43  => ("000101011", "00000000000001010", "00011100101000000"),
    44  => ("000101100", "00000000000001010", "10110111100110000"),
    45  => ("000101101", "00000000000001010", "00000111101110000"),
    46  => ("000101110", "00000000000001010", "00111001110111110"),
    47  => ("000101111", "00000000000001010", "10101011101101100"),
    48  => ("000110000", "00000000000001010", "01000011001111011"),
    49  => ("000110001", "00000000000001010", "11101011001001111"),
    50  => ("000110010", "00000000000001010", "01110110111001110"),
    51  => ("000110011", "00000000000001010", "10101001100100110"),
    52  => ("000110100", "00000000000001010", "01011010001100101"),
    53  => ("000110101", "00000000000001010", "00000000101111000"),
    54  => ("000110110", "00000000000001010", "11111000100000011"),
    55  => ("000110111", "00000000000001010", "10110000111100011"),
    56  => ("000111000", "00000000000001010", "00000100001000011"),
    57  => ("000111001", "00000000000001010", "01111101100010101"),
    58  => ("000111010", "00000000000001010", "11101111111110001"),
    59  => ("000111011", "00000000000001010", "00100001111001001"),
    60  => ("000111100", "00000000000001010", "00011110111101001"),
    61  => ("000111101", "00000000000001010", "01010100001101100"),
    62  => ("000111110", "00000000000001010", "11001010110110010"),
    63  => ("000111111", "00000000000001010", "00110100010001001"),
    64  => ("001000000", "00000000000001010", "00101001100011010"),
    65  => ("001000001", "00000000000001010", "10010001101111000"),
    66  => ("001000010", "00000000000001010", "10010100000010111"),
    67  => ("001000011", "00000000000001010", "10100111000111011"),
    68  => ("001000100", "00000000000001010", "11111011010010110"),
    69  => ("001000101", "00000000000001010", "01110000100100101"),
    70  => ("001000110", "00000000000001010", "00000011011101100"),
    71  => ("001000111", "00000000000001010", "10000100100001101"),
    72  => ("001001000", "00000000000001010", "10101101110101001"),
    73  => ("001001001", "00000000000001010", "01001110011000011"),
    74  => ("001001010", "00000000000001010", "00011110001011100"),
    75  => ("001001011", "00000000000001010", "10110100011010001"),
    76  => ("001001100", "00000000000001010", "11100110110100011"),
    77  => ("001001101", "00000000000001010", "01001010100101011"),
    78  => ("001001110", "00000000000001010", "00001001011011100"),
    79  => ("001001111", "00000000000001010", "11100010101111100"),
    80  => ("001010000", "00000000000001010", "10110101101101011"),
    81  => ("001010001", "00000000000001010", "10101011000000101"),
    82  => ("001010010", "00000000000001010", "01001110001000101"),
    83  => ("001010011", "00000000000001010", "10001011110110110"),
    84  => ("001010100", "00000000000001010", "11110111001100100"),
    85  => ("001010101", "00000000000001010", "10000000100110111"),
    86  => ("001010110", "00000000000001010", "01011100110111111"),
    87  => ("001010111", "00000000000001010", "01101010010010001"),
    88  => ("001011000", "00000000000001010", "00111100100011011"),
    89  => ("001011001", "00000000000001010", "01101001011111110"),
    90  => ("001011010", "00000000000001010", "10100001110100011"),
    91  => ("001011011", "00000000000001010", "00100011011011011"),
    92  => ("001011100", "00000000000001010", "01010100110110011"),
    93  => ("001011101", "00000000000001010", "00100100111000110"),
    94  => ("001011110", "00000000000001010", "01011100001010110"),
    95  => ("001011111", "00000000000001010", "01100000110101000"),
    96  => ("001100000", "00000000000001010", "11111011111011100"),
    97  => ("001100001", "00000000000001010", "10000001001011111"),
    98  => ("001100010", "00000000000001010", "11110110011010000"),
    99  => ("001100011", "00000000000001010", "01000001111101111"),
    100 => ("001100100", "00000000000001010", "10101011011101001"),
    101 => ("001100101", "00000000000001010", "01001001010011010"),
    102 => ("001100110", "00000000000001010", "11010111011111001"),
    103 => ("001100111", "00000000000001010", "01010001010000110"),
    104 => ("001101000", "00000000000001010", "01101111000011100"),
    105 => ("001101001", "00000000000001010", "10011010101010011"),
    106 => ("001101010", "00000000000001010", "00010000010111100"),
    107 => ("001101011", "00000000000001010", "10010011011100100"),
    108 => ("001101100", "00000000000001010", "11100101001100100"),
    109 => ("001101101", "00000000000001010", "01100001001110000"),
    110 => ("001101110", "00000000000001010", "11011011111000101"),
    111 => ("001101111", "00000000000001010", "10000101000001111"),
    112 => ("001110000", "00000000000001010", "01110000111000010"),
    113 => ("001110001", "00000000000001010", "10111111111011111"),
    114 => ("001110010", "00000000000001010", "01001111111100110"),
    115 => ("001110011", "00000000000001010", "10100110111110110"),
    116 => ("001110100", "00000000000001010", "11001111110100110"),
    117 => ("001110101", "00000000000001010", "01010010001100010"),
    118 => ("001110110", "00000000000001010", "10000100011111111"),
    119 => ("001110111", "00000000000001010", "00100110010110111"),
    120 => ("001111000", "00000000000001010", "11110111010101100"),
    121 => ("001111001", "00000000000001010", "00011001001011100"),
    122 => ("001111010", "00000000000001010", "00111110001101100"),
    123 => ("001111011", "00000000000001010", "11010000011010100"),
    124 => ("001111100", "00000000000001010", "11010101011110011"),
    125 => ("001111101", "00000000000001010", "00000011100101010"),
    126 => ("001111110", "00000000000001010", "00110100011111001"),
    127 => ("001111111", "00000000000001010", "01110100010101011"),
    128 => ("010000000", "00000000000001010", "10111101110100001"),
    129 => ("010000001", "00000000000001010", "10100101111110111"),
    130 => ("010000010", "00000000000001010", "10001100100011000"),
    131 => ("010000011", "00000000000001010", "01010110010001010"),
    132 => ("010000100", "00000000000001010", "01010001010000111"),
    133 => ("010000101", "00000000000001010", "11111111001101100"),
    134 => ("010000110", "00000000000001010", "01111000110111011"),
    135 => ("010000111", "00000000000001010", "00000100110101000"),
    136 => ("010001000", "00000000000001010", "01000001010101110"),
    137 => ("010001001", "00000000000001010", "00010010111010011"),
    138 => ("010001010", "00000000000001010", "11100010111111010"),
    139 => ("010001011", "00000000000001010", "01011111110111011"),
    140 => ("010001100", "00000000000001010", "00101100101101100"),
    141 => ("010001101", "00000000000001010", "10000110101001100"),
    142 => ("010001110", "00000000000001010", "01111111110111101"),
    143 => ("010001111", "00000000000001010", "01111111111011001"),
    144 => ("010010000", "00000000000001010", "00010100001001001"),
    145 => ("010010001", "00000000000001010", "00100000001011110"),
    146 => ("010010010", "00000000000001010", "10101011010010101"),
    147 => ("010010011", "00000000000001010", "10000111111010100"),
    148 => ("010010100", "00000000000001010", "11010001011111100"),
    149 => ("010010101", "00000000000001010", "10011100101100101"),
    150 => ("010010110", "00000000000001010", "10101010001100100"),
    151 => ("010010111", "00000000000001010", "11101111011101100"),
    152 => ("010011000", "00000000000001010", "01001101001010011"),
    153 => ("010011001", "00000000000001010", "10001111011000010"),
    154 => ("010011010", "00000000000001010", "10001000011001101"),
    155 => ("010011011", "00000000000001010", "11001011011101000"),
    156 => ("010011100", "00000000000001010", "01010001100001000"),
    157 => ("010011101", "00000000000001010", "01100001111110010"),
    158 => ("010011110", "00000000000001010", "11111101111110111"),
    159 => ("010011111", "00000000000001010", "01011101001101111"),
    160 => ("010100000", "00000000000001010", "10100110001110110"),
    161 => ("010100001", "00000000000001010", "11101101011001001"),
    162 => ("010100010", "00000000000001010", "01100100001000010"),
    163 => ("010100011", "00000000000001010", "10000111111110111"),
    164 => ("010100100", "00000000000001010", "01111101100000000"),
    165 => ("010100101", "00000000000001010", "00110011111110011"),
    166 => ("010100110", "00000000000001010", "00110111011010000"),
    167 => ("010100111", "00000000000001010", "01010001110001110"),
    168 => ("010101000", "00000000000001010", "10000011001001010"),
    169 => ("010101001", "00000000000001010", "00000011000101110"),
    170 => ("010101010", "00000000000001010", "00111011010111000"),
    171 => ("010101011", "00000000000001010", "00111011111100100"),
    172 => ("010101100", "00000000000001010", "00001101000010011"),
    173 => ("010101101", "00000000000001010", "10100110001111000"),
    174 => ("010101110", "00000000000001010", "01010011010110010"),
    175 => ("010101111", "00000000000001010", "11011110010001110"),
    176 => ("010110000", "00000000000001010", "10100101100000110"),
    177 => ("010110001", "00000000000001010", "11011001100010100"),
    178 => ("010110010", "00000000000001010", "10111010000000010"),
    179 => ("010110011", "00000000000001010", "10011010110010001"),
    180 => ("010110100", "00000000000001010", "10001100110010110"),
    181 => ("010110101", "00000000000001010", "01100111000100100"),
    182 => ("010110110", "00000000000001010", "11000111010100001"),
    183 => ("010110111", "00000000000001010", "01110110000110101"),
    184 => ("010111000", "00000000000001010", "11101000010001110"),
    185 => ("010111001", "00000000000001010", "01111100100001100"),
    186 => ("010111010", "00000000000001010", "10000010101101101"),
    187 => ("010111011", "00000000000001010", "00010110011010000"),
    188 => ("010111100", "00000000000001010", "10110010101111111"),
    189 => ("010111101", "00000000000001010", "01001100111011001"),
    190 => ("010111110", "00000000000001010", "00100010100001100"),
    191 => ("010111111", "00000000000001010", "10110100011110011"),
    192 => ("011000000", "00000000000001010", "11100010001101111"),
    193 => ("011000001", "00000000000001010", "01000101010011111"),
    194 => ("011000010", "00000000000001010", "10101101110010101"),
    195 => ("011000011", "00000000000001010", "00101010001010110"),
    196 => ("011000100", "00000000000001010", "10111001001011110"),
    197 => ("011000101", "00000000000001010", "01011110101100000"),
    198 => ("011000110", "00000000000001010", "01011001101100000"),
    199 => ("011000111", "00000000000001010", "00001111010001100"),
    200 => ("011001000", "00000000000001010", "11001001111000100"),
    201 => ("011001001", "00000000000001010", "01100111101011011"),
    202 => ("011001010", "00000000000001010", "11010000010010000"),
    203 => ("011001011", "00000000000001010", "00001001000010011"),
    204 => ("011001100", "00000000000001010", "11100010101011100"),
    205 => ("011001101", "00000000000001010", "11001001010010111"),
    206 => ("011001110", "00000000000001010", "01111110001101001"),
    207 => ("011001111", "00000000000001010", "10011100000001001"),
    208 => ("011010000", "00000000000001010", "01011101101100010"),
    209 => ("011010001", "00000000000001010", "10000111111110000"),
    210 => ("011010010", "00000000000001010", "01110001101100111"),
    211 => ("011010011", "00000000000001010", "00000101110000001"),
    212 => ("011010100", "00000000000001010", "01001010000100110"),
    213 => ("011010101", "00000000000001010", "00101001011110101"),
    214 => ("011010110", "00000000000001010", "01110110010111010"),
    215 => ("011010111", "00000000000001010", "11000011110000101"),
    216 => ("011011000", "00000000000001010", "10100000000000011"),
    217 => ("011011001", "00000000000001010", "10010010101000110"),
    218 => ("011011010", "00000000000001010", "10110000100100101"),
    219 => ("011011011", "00000000000001010", "00001001010010111"),
    220 => ("011011100", "00000000000001010", "11001101101001101"),
    221 => ("011011101", "00000000000001010", "11111001111101010"),
    222 => ("011011110", "00000000000001010", "00011110001011101"),
    223 => ("011011111", "00000000000001010", "11101101010000001"),
    224 => ("011100000", "00000000000001010", "00000001010101100"),
    225 => ("011100001", "00000000000001010", "00000000100101110"),
    226 => ("011100010", "00000000000001010", "01101111001100001"),
    227 => ("011100011", "00000000000001010", "10111011101111011"),
    228 => ("011100100", "00000000000001010", "01011110100000110"),
    229 => ("011100101", "00000000000001010", "11111110011000100"),
    230 => ("011100110", "00000000000001010", "10101111110111010"),
    231 => ("011100111", "00000000000001010", "00100110101100010"),
    232 => ("011101000", "00000000000001010", "01110111110011010"),
    233 => ("011101001", "00000000000001010", "01101110010011111"),
    234 => ("011101010", "00000000000001010", "10010100110111101"),
    235 => ("011101011", "00000000000001010", "11001100001111000"),
    236 => ("011101100", "00000000000001010", "11111010011110011"),
    237 => ("011101101", "00000000000001010", "10111011010011111"),
    238 => ("011101110", "00000000000001010", "00111101111001010"),
    239 => ("011101111", "00000000000001010", "10010101011111101"),
    240 => ("011110000", "00000000000001010", "00001100011011010"),
    241 => ("011110001", "00000000000001010", "10000101010010011"),
    242 => ("011110010", "00000000000001010", "00101110000110101"),
    243 => ("011110011", "00000000000001010", "00101001000011000"),
    244 => ("011110100", "00000000000001010", "11010100000111100"),
    245 => ("011110101", "00000000000001010", "00110100101001011"),
    246 => ("011110110", "00000000000001010", "01011001111011100"),
    247 => ("011110111", "00000000000001010", "11100000010111100"),
    248 => ("011111000", "00000000000001010", "11101100110100010"),
    249 => ("011111001", "00000000000001010", "10110001001101111"),
    250 => ("011111010", "00000000000001010", "11111110101010111"),
    251 => ("011111011", "00000000000001010", "10101011110010010"),
    252 => ("011111100", "00000000000001010", "01110101111010000"),
    253 => ("011111101", "00000000000001010", "01101010010011100"),
    254 => ("011111110", "00000000000001010", "01101111011011011"),
    255 => ("011111111", "00000000000001010", "10011111010100011")
  );

end package;
